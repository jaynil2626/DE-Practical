<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>303.251,5.40273,425.789,-55.1656</PageViewport>
<gate>
<ID>193</ID>
<type>AA_TOGGLE</type>
<position>342,-8</position>
<output>
<ID>OUT_0</ID>102 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>194</ID>
<type>AA_TOGGLE</type>
<position>347,-8</position>
<output>
<ID>OUT_0</ID>100 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>195</ID>
<type>AA_TOGGLE</type>
<position>352,-8</position>
<output>
<ID>OUT_0</ID>99 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>2</ID>
<type>AA_MUX_2x1</type>
<position>22,-13.5</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>4 </output>
<input>
<ID>SEL_0</ID>3 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>196</ID>
<type>AA_TOGGLE</type>
<position>357,-8</position>
<output>
<ID>OUT_0</ID>98 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>197</ID>
<type>AA_TOGGLE</type>
<position>362,-8</position>
<output>
<ID>OUT_0</ID>97 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>15.5,-12</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>199</ID>
<type>AE_OR4</type>
<position>371,-16</position>
<input>
<ID>IN_0</ID>100 </input>
<input>
<ID>IN_1</ID>99 </input>
<input>
<ID>IN_2</ID>98 </input>
<input>
<ID>IN_3</ID>97 </input>
<output>
<ID>OUT</ID>104 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>15.5,-15</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>200</ID>
<type>AE_OR4</type>
<position>371,-28</position>
<input>
<ID>IN_0</ID>101 </input>
<input>
<ID>IN_1</ID>102 </input>
<input>
<ID>IN_2</ID>98 </input>
<input>
<ID>IN_3</ID>97 </input>
<output>
<ID>OUT</ID>105 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>201</ID>
<type>AE_OR4</type>
<position>371,-40</position>
<input>
<ID>IN_0</ID>103 </input>
<input>
<ID>IN_1</ID>102 </input>
<input>
<ID>IN_2</ID>99 </input>
<input>
<ID>IN_3</ID>97 </input>
<output>
<ID>OUT</ID>106 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>22,-8</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>203</ID>
<type>GA_LED</type>
<position>379,-16</position>
<input>
<ID>N_in0</ID>104 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>GA_LED</type>
<position>26.5,-13.5</position>
<input>
<ID>N_in0</ID>4 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>205</ID>
<type>GA_LED</type>
<position>379,-28</position>
<input>
<ID>N_in0</ID>105 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>AA_LABEL</type>
<position>22,-1.5</position>
<gparam>LABEL_TEXT 2x1 MUX</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>207</ID>
<type>GA_LED</type>
<position>379,-40</position>
<input>
<ID>N_in0</ID>106 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>AE_MUX_4x1</type>
<position>49.5,-14</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>7 </input>
<input>
<ID>IN_2</ID>6 </input>
<input>
<ID>IN_3</ID>5 </input>
<output>
<ID>OUT</ID>11 </output>
<input>
<ID>SEL_0</ID>10 </input>
<input>
<ID>SEL_1</ID>9 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>208</ID>
<type>AA_LABEL</type>
<position>327,-4</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>209</ID>
<type>AA_LABEL</type>
<position>332,-4</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>AA_TOGGLE</type>
<position>43.5,-11</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>210</ID>
<type>AA_LABEL</type>
<position>337,-4</position>
<gparam>LABEL_TEXT D2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>211</ID>
<type>AA_LABEL</type>
<position>342,-4</position>
<gparam>LABEL_TEXT D3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>AA_TOGGLE</type>
<position>43.5,-13</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>212</ID>
<type>AA_LABEL</type>
<position>346.5,-4</position>
<gparam>LABEL_TEXT D4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>213</ID>
<type>AA_LABEL</type>
<position>352,-4</position>
<gparam>LABEL_TEXT D5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>AA_TOGGLE</type>
<position>43.5,-15</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>214</ID>
<type>AA_LABEL</type>
<position>357,-4</position>
<gparam>LABEL_TEXT D6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>215</ID>
<type>AA_LABEL</type>
<position>362,-4</position>
<gparam>LABEL_TEXT D7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>AA_TOGGLE</type>
<position>43.5,-17</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>216</ID>
<type>AA_LABEL</type>
<position>383,-15.5</position>
<gparam>LABEL_TEXT S2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>217</ID>
<type>AA_LABEL</type>
<position>383,-27.5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>AA_TOGGLE</type>
<position>48.5,-6</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>218</ID>
<type>AA_LABEL</type>
<position>383,-39.5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>219</ID>
<type>AA_LABEL</type>
<position>348,-0.5</position>
<gparam>LABEL_TEXT 8x3 Encoder (octal to binary)</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>AA_TOGGLE</type>
<position>51.5,-6</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>28</ID>
<type>GA_LED</type>
<position>56,-14</position>
<input>
<ID>N_in0</ID>11 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>29</ID>
<type>AA_LABEL</type>
<position>50,-1.5</position>
<gparam>LABEL_TEXT 4x1 MUX</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>31</ID>
<type>AI_MUX_8x1</type>
<position>82,-16</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>18 </input>
<input>
<ID>IN_2</ID>17 </input>
<input>
<ID>IN_3</ID>16 </input>
<input>
<ID>IN_4</ID>15 </input>
<input>
<ID>IN_5</ID>14 </input>
<input>
<ID>IN_6</ID>13 </input>
<input>
<ID>IN_7</ID>12 </input>
<output>
<ID>OUT</ID>23 </output>
<input>
<ID>SEL_0</ID>22 </input>
<input>
<ID>SEL_1</ID>21 </input>
<input>
<ID>SEL_2</ID>20 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>33</ID>
<type>AA_TOGGLE</type>
<position>71,-9.5</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>35</ID>
<type>AA_TOGGLE</type>
<position>71,-11.5</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>37</ID>
<type>AA_TOGGLE</type>
<position>71,-13.5</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>39</ID>
<type>AA_TOGGLE</type>
<position>71,-15.5</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>41</ID>
<type>AA_TOGGLE</type>
<position>71,-17.5</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>43</ID>
<type>AA_TOGGLE</type>
<position>71,-19.5</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>45</ID>
<type>AA_TOGGLE</type>
<position>71,-21.5</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>47</ID>
<type>AA_TOGGLE</type>
<position>71,-23.5</position>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>49</ID>
<type>AA_TOGGLE</type>
<position>79,-6</position>
<output>
<ID>OUT_0</ID>20 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>51</ID>
<type>AA_TOGGLE</type>
<position>82,-6</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>53</ID>
<type>AA_TOGGLE</type>
<position>85,-6</position>
<output>
<ID>OUT_0</ID>22 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>55</ID>
<type>GA_LED</type>
<position>87,-16</position>
<input>
<ID>N_in0</ID>23 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>56</ID>
<type>AA_LABEL</type>
<position>81.5,-1.5</position>
<gparam>LABEL_TEXT 8x1 MUX</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>61</ID>
<type>AA_MUX_2x1</type>
<position>119.5,-13.5</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>44 </output>
<input>
<ID>SEL_0</ID>26 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>62</ID>
<type>AA_TOGGLE</type>
<position>113,-12</position>
<output>
<ID>OUT_0</ID>24 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>63</ID>
<type>AA_TOGGLE</type>
<position>113,-15</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>64</ID>
<type>AA_TOGGLE</type>
<position>119.5,-8</position>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>66</ID>
<type>AA_MUX_2x1</type>
<position>119.5,-23.5</position>
<input>
<ID>IN_0</ID>29 </input>
<input>
<ID>IN_1</ID>28 </input>
<output>
<ID>OUT</ID>45 </output>
<input>
<ID>SEL_0</ID>26 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>67</ID>
<type>AA_TOGGLE</type>
<position>113,-22</position>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>68</ID>
<type>AA_TOGGLE</type>
<position>113,-25</position>
<output>
<ID>OUT_0</ID>29 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>71</ID>
<type>AA_MUX_2x1</type>
<position>119.5,-33.5</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>50 </output>
<input>
<ID>SEL_0</ID>26 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>72</ID>
<type>AA_TOGGLE</type>
<position>113,-32</position>
<output>
<ID>OUT_0</ID>32 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>73</ID>
<type>AA_TOGGLE</type>
<position>113,-35</position>
<output>
<ID>OUT_0</ID>33 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>76</ID>
<type>AA_MUX_2x1</type>
<position>119.5,-43.5</position>
<input>
<ID>IN_0</ID>37 </input>
<input>
<ID>IN_1</ID>36 </input>
<output>
<ID>OUT</ID>51 </output>
<input>
<ID>SEL_0</ID>26 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>77</ID>
<type>AA_TOGGLE</type>
<position>113,-42</position>
<output>
<ID>OUT_0</ID>36 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>78</ID>
<type>AA_TOGGLE</type>
<position>113,-45</position>
<output>
<ID>OUT_0</ID>37 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>81</ID>
<type>AA_MUX_2x1</type>
<position>131,-22.5</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>IN_1</ID>44 </input>
<output>
<ID>OUT</ID>57 </output>
<input>
<ID>SEL_0</ID>42 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>84</ID>
<type>AA_TOGGLE</type>
<position>131,-8</position>
<output>
<ID>OUT_0</ID>42 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>86</ID>
<type>AA_MUX_2x1</type>
<position>131,-34.5</position>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>50 </input>
<output>
<ID>OUT</ID>56 </output>
<input>
<ID>SEL_0</ID>42 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>93</ID>
<type>AA_MUX_2x1</type>
<position>143,-27.5</position>
<input>
<ID>IN_0</ID>56 </input>
<input>
<ID>IN_1</ID>57 </input>
<output>
<ID>OUT</ID>55 </output>
<input>
<ID>SEL_0</ID>54 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>96</ID>
<type>AA_TOGGLE</type>
<position>143,-8</position>
<output>
<ID>OUT_0</ID>54 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>97</ID>
<type>GA_LED</type>
<position>147.5,-27.5</position>
<input>
<ID>N_in0</ID>55 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>98</ID>
<type>AA_LABEL</type>
<position>130,-1.5</position>
<gparam>LABEL_TEXT 8x1 using 2x1 MUX</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>100</ID>
<type>AA_LABEL</type>
<position>109,-11.5</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>101</ID>
<type>AA_LABEL</type>
<position>109,-15</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>102</ID>
<type>AA_LABEL</type>
<position>109,-21.5</position>
<gparam>LABEL_TEXT D2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>103</ID>
<type>AA_LABEL</type>
<position>109,-24.5</position>
<gparam>LABEL_TEXT D3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>104</ID>
<type>AA_LABEL</type>
<position>109,-32</position>
<gparam>LABEL_TEXT D4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>105</ID>
<type>AA_LABEL</type>
<position>109,-35</position>
<gparam>LABEL_TEXT D5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>106</ID>
<type>AA_LABEL</type>
<position>109,-42</position>
<gparam>LABEL_TEXT D6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>107</ID>
<type>AA_LABEL</type>
<position>109,-45</position>
<gparam>LABEL_TEXT D7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>108</ID>
<type>AA_LABEL</type>
<position>143,-5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>109</ID>
<type>AA_LABEL</type>
<position>131,-5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>110</ID>
<type>AA_LABEL</type>
<position>119.5,-5</position>
<gparam>LABEL_TEXT S2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>115</ID>
<type>AA_TOGGLE</type>
<position>169.5,-8</position>
<output>
<ID>OUT_0</ID>58 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>117</ID>
<type>AA_TOGGLE</type>
<position>178,-8</position>
<output>
<ID>OUT_0</ID>61 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>119</ID>
<type>AA_TOGGLE</type>
<position>185.5,-8</position>
<output>
<ID>OUT_0</ID>59 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>123</ID>
<type>AA_AND3</type>
<position>202,-15</position>
<input>
<ID>IN_0</ID>59 </input>
<input>
<ID>IN_1</ID>67 </input>
<input>
<ID>IN_2</ID>60 </input>
<output>
<ID>OUT</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>125</ID>
<type>AA_AND3</type>
<position>202,-24</position>
<input>
<ID>IN_0</ID>59 </input>
<input>
<ID>IN_1</ID>60 </input>
<input>
<ID>IN_2</ID>61 </input>
<output>
<ID>OUT</ID>64 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>127</ID>
<type>AA_AND3</type>
<position>202,-32</position>
<input>
<ID>IN_0</ID>59 </input>
<input>
<ID>IN_1</ID>58 </input>
<input>
<ID>IN_2</ID>67 </input>
<output>
<ID>OUT</ID>65 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>129</ID>
<type>AA_AND3</type>
<position>202,-40</position>
<input>
<ID>IN_0</ID>59 </input>
<input>
<ID>IN_1</ID>58 </input>
<input>
<ID>IN_2</ID>61 </input>
<output>
<ID>OUT</ID>66 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>133</ID>
<type>AE_SMALL_INVERTER</type>
<position>171.5,-11</position>
<input>
<ID>IN_0</ID>58 </input>
<output>
<ID>OUT_0</ID>60 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>135</ID>
<type>AE_SMALL_INVERTER</type>
<position>180,-11</position>
<input>
<ID>IN_0</ID>61 </input>
<output>
<ID>OUT_0</ID>67 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>139</ID>
<type>GA_LED</type>
<position>210.5,-15</position>
<input>
<ID>N_in0</ID>63 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>141</ID>
<type>GA_LED</type>
<position>210.5,-24</position>
<input>
<ID>N_in0</ID>64 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>143</ID>
<type>GA_LED</type>
<position>210.5,-32</position>
<input>
<ID>N_in0</ID>65 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>145</ID>
<type>GA_LED</type>
<position>210.5,-40</position>
<input>
<ID>N_in0</ID>66 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>147</ID>
<type>AA_LABEL</type>
<position>189.5,-1.5</position>
<gparam>LABEL_TEXT 1x4 Demux</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>148</ID>
<type>AA_LABEL</type>
<position>178,-5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>149</ID>
<type>AA_LABEL</type>
<position>169.5,-5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>150</ID>
<type>AA_LABEL</type>
<position>185.5,-5</position>
<gparam>LABEL_TEXT Din</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>151</ID>
<type>AA_TOGGLE</type>
<position>258,-8</position>
<output>
<ID>OUT_0</ID>68 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>152</ID>
<type>AA_TOGGLE</type>
<position>266.5,-8</position>
<output>
<ID>OUT_0</ID>71 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>153</ID>
<type>AA_TOGGLE</type>
<position>274,-8</position>
<output>
<ID>OUT_0</ID>86 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>158</ID>
<type>AE_SMALL_INVERTER</type>
<position>260,-11</position>
<input>
<ID>IN_0</ID>68 </input>
<output>
<ID>OUT_0</ID>84 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>159</ID>
<type>AE_SMALL_INVERTER</type>
<position>268.5,-11</position>
<input>
<ID>IN_0</ID>71 </input>
<output>
<ID>OUT_0</ID>85 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>160</ID>
<type>GA_LED</type>
<position>293.5,-17</position>
<input>
<ID>N_in0</ID>77 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>161</ID>
<type>GA_LED</type>
<position>293.5,-27</position>
<input>
<ID>N_in0</ID>78 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>162</ID>
<type>GA_LED</type>
<position>293.5,-37</position>
<input>
<ID>N_in0</ID>79 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>163</ID>
<type>GA_LED</type>
<position>293.5,-47</position>
<input>
<ID>N_in0</ID>80 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>164</ID>
<type>AA_LABEL</type>
<position>266.5,-5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>165</ID>
<type>AA_LABEL</type>
<position>258,-5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>166</ID>
<type>AA_LABEL</type>
<position>274,-5</position>
<gparam>LABEL_TEXT Din</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>168</ID>
<type>AA_AND4</type>
<position>287,-17</position>
<input>
<ID>IN_0</ID>83 </input>
<input>
<ID>IN_1</ID>84 </input>
<input>
<ID>IN_2</ID>85 </input>
<input>
<ID>IN_3</ID>86 </input>
<output>
<ID>OUT</ID>77 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>169</ID>
<type>AA_AND4</type>
<position>287,-27</position>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>84 </input>
<input>
<ID>IN_2</ID>85 </input>
<input>
<ID>IN_3</ID>86 </input>
<output>
<ID>OUT</ID>78 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>170</ID>
<type>AA_AND4</type>
<position>287,-37</position>
<input>
<ID>IN_0</ID>83 </input>
<input>
<ID>IN_1</ID>68 </input>
<input>
<ID>IN_2</ID>85 </input>
<input>
<ID>IN_3</ID>86 </input>
<output>
<ID>OUT</ID>79 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>171</ID>
<type>AA_AND4</type>
<position>287,-47</position>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>68 </input>
<input>
<ID>IN_2</ID>85 </input>
<input>
<ID>IN_3</ID>86 </input>
<output>
<ID>OUT</ID>80 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>172</ID>
<type>AA_TOGGLE</type>
<position>249.5,-8</position>
<output>
<ID>OUT_0</ID>81 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>173</ID>
<type>AE_SMALL_INVERTER</type>
<position>251.5,-11</position>
<input>
<ID>IN_0</ID>81 </input>
<output>
<ID>OUT_0</ID>83 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>176</ID>
<type>AA_LABEL</type>
<position>249.5,-5</position>
<gparam>LABEL_TEXT S2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>178</ID>
<type>GA_LED</type>
<position>293.5,-57</position>
<input>
<ID>N_in0</ID>88 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>179</ID>
<type>GA_LED</type>
<position>293.5,-67</position>
<input>
<ID>N_in0</ID>89 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>180</ID>
<type>GA_LED</type>
<position>293.5,-77</position>
<input>
<ID>N_in0</ID>90 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>181</ID>
<type>GA_LED</type>
<position>293.5,-87</position>
<input>
<ID>N_in0</ID>91 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>182</ID>
<type>AA_AND4</type>
<position>287,-57</position>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>84 </input>
<input>
<ID>IN_2</ID>83 </input>
<input>
<ID>IN_3</ID>86 </input>
<output>
<ID>OUT</ID>88 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>183</ID>
<type>AA_AND4</type>
<position>287,-67</position>
<input>
<ID>IN_0</ID>83 </input>
<input>
<ID>IN_1</ID>68 </input>
<input>
<ID>IN_2</ID>85 </input>
<input>
<ID>IN_3</ID>86 </input>
<output>
<ID>OUT</ID>89 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>184</ID>
<type>AA_AND4</type>
<position>287,-77</position>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>68 </input>
<input>
<ID>IN_2</ID>83 </input>
<input>
<ID>IN_3</ID>86 </input>
<output>
<ID>OUT</ID>90 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>185</ID>
<type>AA_AND4</type>
<position>287,-87</position>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>68 </input>
<input>
<ID>IN_2</ID>71 </input>
<input>
<ID>IN_3</ID>86 </input>
<output>
<ID>OUT</ID>91 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>186</ID>
<type>AA_LABEL</type>
<position>272,-0.5</position>
<gparam>LABEL_TEXT 1x8 Demux</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>188</ID>
<type>AA_TOGGLE</type>
<position>327,-8</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>190</ID>
<type>AA_TOGGLE</type>
<position>332,-8</position>
<output>
<ID>OUT_0</ID>103 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>192</ID>
<type>AA_TOGGLE</type>
<position>337,-8</position>
<output>
<ID>OUT_0</ID>101 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,-12.5,20,-12</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,-12,20,-12</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>20 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,-15,20,-14.5</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,-15,20,-15</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>20 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-11,22,-10</points>
<connection>
<GID>2</GID>
<name>SEL_0</name></connection>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24,-13.5,25.5,-13.5</points>
<connection>
<GID>10</GID>
<name>N_in0</name></connection>
<connection>
<GID>2</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-11,46.5,-11</points>
<connection>
<GID>14</GID>
<name>IN_3</name></connection>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-13,46.5,-13</points>
<connection>
<GID>14</GID>
<name>IN_2</name></connection>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-15,46.5,-15</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>46.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>46.5,-15,46.5,-15</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>-15 1</intersection></vsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-17,46.5,-17</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<intersection>46.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>46.5,-17,46.5,-17</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>-17 1</intersection></vsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-9,49.5,-8.5</points>
<connection>
<GID>14</GID>
<name>SEL_1</name></connection>
<intersection>-8.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>48.5,-8.5,48.5,-8</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>-8.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-8.5,49.5,-8.5</points>
<intersection>48.5 1</intersection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-9,50.5,-8.5</points>
<connection>
<GID>14</GID>
<name>SEL_0</name></connection>
<intersection>-8.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>51.5,-8.5,51.5,-8</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>-8.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>50.5,-8.5,51.5,-8.5</points>
<intersection>50.5 0</intersection>
<intersection>51.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>52.5,-14,55,-14</points>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<connection>
<GID>28</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78,-12.5,78,-9.5</points>
<intersection>-12.5 1</intersection>
<intersection>-9.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>78,-12.5,79,-12.5</points>
<connection>
<GID>31</GID>
<name>IN_7</name></connection>
<intersection>78 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>73,-9.5,78,-9.5</points>
<connection>
<GID>33</GID>
<name>OUT_0</name></connection>
<intersection>78 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>77,-13.5,79,-13.5</points>
<connection>
<GID>31</GID>
<name>IN_6</name></connection>
<intersection>77 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>77,-13.5,77,-11.5</points>
<intersection>-13.5 1</intersection>
<intersection>-11.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>73,-11.5,77,-11.5</points>
<connection>
<GID>35</GID>
<name>OUT_0</name></connection>
<intersection>77 4</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-14.5,76,-13.5</points>
<intersection>-14.5 1</intersection>
<intersection>-13.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76,-14.5,79,-14.5</points>
<connection>
<GID>31</GID>
<name>IN_5</name></connection>
<intersection>76 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>73,-13.5,76,-13.5</points>
<connection>
<GID>37</GID>
<name>OUT_0</name></connection>
<intersection>76 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-15.5,79,-15.5</points>
<connection>
<GID>39</GID>
<name>OUT_0</name></connection>
<connection>
<GID>31</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-17.5,76,-16.5</points>
<intersection>-17.5 2</intersection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76,-16.5,79,-16.5</points>
<connection>
<GID>31</GID>
<name>IN_3</name></connection>
<intersection>76 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>73,-17.5,76,-17.5</points>
<connection>
<GID>41</GID>
<name>OUT_0</name></connection>
<intersection>76 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77,-19.5,77,-17.5</points>
<intersection>-19.5 2</intersection>
<intersection>-17.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77,-17.5,79,-17.5</points>
<connection>
<GID>31</GID>
<name>IN_2</name></connection>
<intersection>77 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>73,-19.5,77,-19.5</points>
<connection>
<GID>43</GID>
<name>OUT_0</name></connection>
<intersection>77 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78,-21.5,78,-18.5</points>
<intersection>-21.5 2</intersection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>78,-18.5,79,-18.5</points>
<connection>
<GID>31</GID>
<name>IN_1</name></connection>
<intersection>78 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>73,-21.5,78,-21.5</points>
<connection>
<GID>45</GID>
<name>OUT_0</name></connection>
<intersection>78 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79,-23.5,79,-19.5</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>-23.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>73,-23.5,79,-23.5</points>
<connection>
<GID>47</GID>
<name>OUT_0</name></connection>
<intersection>79 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,-10.5,81,-8.5</points>
<connection>
<GID>31</GID>
<name>SEL_2</name></connection>
<intersection>-8.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>79,-8.5,79,-8</points>
<connection>
<GID>49</GID>
<name>OUT_0</name></connection>
<intersection>-8.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>79,-8.5,81,-8.5</points>
<intersection>79 1</intersection>
<intersection>81 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>6</ID>
<points>82,-10.5,82,-8</points>
<connection>
<GID>51</GID>
<name>OUT_0</name></connection>
<intersection>-10.5 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>82,-10.5,82,-10.5</points>
<connection>
<GID>31</GID>
<name>SEL_1</name></connection>
<intersection>82 6</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83,-10.5,83,-8.5</points>
<connection>
<GID>31</GID>
<name>SEL_0</name></connection>
<intersection>-8.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>85,-8.5,85,-8</points>
<connection>
<GID>53</GID>
<name>OUT_0</name></connection>
<intersection>-8.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>83,-8.5,85,-8.5</points>
<intersection>83 0</intersection>
<intersection>85 1</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>85,-16,86,-16</points>
<connection>
<GID>55</GID>
<name>N_in0</name></connection>
<connection>
<GID>31</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,-12.5,117.5,-12</points>
<connection>
<GID>61</GID>
<name>IN_1</name></connection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115,-12,117.5,-12</points>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection>
<intersection>117.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,-15,117.5,-14.5</points>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115,-15,117.5,-15</points>
<connection>
<GID>63</GID>
<name>OUT_0</name></connection>
<intersection>117.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119.5,-41,119.5,-10</points>
<connection>
<GID>71</GID>
<name>SEL_0</name></connection>
<connection>
<GID>64</GID>
<name>OUT_0</name></connection>
<connection>
<GID>61</GID>
<name>SEL_0</name></connection>
<connection>
<GID>66</GID>
<name>SEL_0</name></connection>
<connection>
<GID>76</GID>
<name>SEL_0</name></connection></vsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,-22.5,117.5,-22</points>
<connection>
<GID>66</GID>
<name>IN_1</name></connection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115,-22,117.5,-22</points>
<connection>
<GID>67</GID>
<name>OUT_0</name></connection>
<intersection>117.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,-25,117.5,-24.5</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>-25 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115,-25,117.5,-25</points>
<connection>
<GID>68</GID>
<name>OUT_0</name></connection>
<intersection>117.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,-32.5,117.5,-32</points>
<connection>
<GID>71</GID>
<name>IN_1</name></connection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115,-32,117.5,-32</points>
<connection>
<GID>72</GID>
<name>OUT_0</name></connection>
<intersection>117.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,-35,117.5,-34.5</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115,-35,117.5,-35</points>
<connection>
<GID>73</GID>
<name>OUT_0</name></connection>
<intersection>117.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,-42.5,117.5,-42</points>
<connection>
<GID>76</GID>
<name>IN_1</name></connection>
<intersection>-42 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115,-42,117.5,-42</points>
<connection>
<GID>77</GID>
<name>OUT_0</name></connection>
<intersection>117.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,-45,117.5,-44.5</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>-45 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115,-45,117.5,-45</points>
<connection>
<GID>78</GID>
<name>OUT_0</name></connection>
<intersection>117.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131,-32,131,-10</points>
<connection>
<GID>84</GID>
<name>OUT_0</name></connection>
<connection>
<GID>81</GID>
<name>SEL_0</name></connection>
<connection>
<GID>86</GID>
<name>SEL_0</name></connection></vsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,-21.5,125,-13.5</points>
<intersection>-21.5 2</intersection>
<intersection>-13.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121.5,-13.5,125,-13.5</points>
<connection>
<GID>61</GID>
<name>OUT</name></connection>
<intersection>125 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>125,-21.5,129,-21.5</points>
<connection>
<GID>81</GID>
<name>IN_1</name></connection>
<intersection>125 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>121.5,-23.5,129,-23.5</points>
<connection>
<GID>81</GID>
<name>IN_0</name></connection>
<connection>
<GID>66</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>121.5,-33.5,129,-33.5</points>
<connection>
<GID>86</GID>
<name>IN_1</name></connection>
<connection>
<GID>71</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,-43.5,125,-35.5</points>
<intersection>-43.5 1</intersection>
<intersection>-35.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121.5,-43.5,125,-43.5</points>
<connection>
<GID>76</GID>
<name>OUT</name></connection>
<intersection>125 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>125,-35.5,129,-35.5</points>
<connection>
<GID>86</GID>
<name>IN_0</name></connection>
<intersection>125 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>143,-25,143,-10</points>
<connection>
<GID>93</GID>
<name>SEL_0</name></connection>
<connection>
<GID>96</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>145,-27.5,146.5,-27.5</points>
<connection>
<GID>97</GID>
<name>N_in0</name></connection>
<connection>
<GID>93</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137,-34.5,137,-28.5</points>
<intersection>-34.5 2</intersection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>137,-28.5,141,-28.5</points>
<connection>
<GID>93</GID>
<name>IN_0</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>133,-34.5,137,-34.5</points>
<connection>
<GID>86</GID>
<name>OUT</name></connection>
<intersection>137 0</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137,-26.5,137,-22.5</points>
<intersection>-26.5 1</intersection>
<intersection>-22.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>137,-26.5,141,-26.5</points>
<connection>
<GID>93</GID>
<name>IN_1</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>133,-22.5,137,-22.5</points>
<connection>
<GID>81</GID>
<name>OUT</name></connection>
<intersection>137 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169.5,-40,169.5,-10</points>
<connection>
<GID>133</GID>
<name>IN_0</name></connection>
<connection>
<GID>115</GID>
<name>OUT_0</name></connection>
<intersection>-40 5</intersection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>169.5,-32,199,-32</points>
<connection>
<GID>127</GID>
<name>IN_1</name></connection>
<intersection>169.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>169.5,-40,199,-40</points>
<connection>
<GID>129</GID>
<name>IN_1</name></connection>
<intersection>169.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185.5,-38,185.5,-10</points>
<connection>
<GID>119</GID>
<name>OUT_0</name></connection>
<intersection>-38 3</intersection>
<intersection>-30 1</intersection>
<intersection>-22 6</intersection>
<intersection>-13 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>185.5,-30,199,-30</points>
<connection>
<GID>127</GID>
<name>IN_0</name></connection>
<intersection>185.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>185.5,-38,199,-38</points>
<connection>
<GID>129</GID>
<name>IN_0</name></connection>
<intersection>185.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>185.5,-13,199,-13</points>
<connection>
<GID>123</GID>
<name>IN_0</name></connection>
<intersection>185.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>185.5,-22,199,-22</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<intersection>185.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>173.5,-24,173.5,-11</points>
<connection>
<GID>133</GID>
<name>OUT_0</name></connection>
<intersection>-24 2</intersection>
<intersection>-17 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>173.5,-24,199,-24</points>
<connection>
<GID>125</GID>
<name>IN_1</name></connection>
<intersection>173.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>173.5,-17,199,-17</points>
<connection>
<GID>123</GID>
<name>IN_2</name></connection>
<intersection>173.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>178,-42,178,-10</points>
<connection>
<GID>117</GID>
<name>OUT_0</name></connection>
<intersection>-42 1</intersection>
<intersection>-26 4</intersection>
<intersection>-11 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>178,-42,199,-42</points>
<connection>
<GID>129</GID>
<name>IN_2</name></connection>
<intersection>178 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>178,-26,199,-26</points>
<connection>
<GID>125</GID>
<name>IN_2</name></connection>
<intersection>178 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>178,-11,178,-11</points>
<connection>
<GID>135</GID>
<name>IN_0</name></connection>
<intersection>178 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>205,-15,209.5,-15</points>
<connection>
<GID>139</GID>
<name>N_in0</name></connection>
<connection>
<GID>123</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>205,-24,209.5,-24</points>
<connection>
<GID>141</GID>
<name>N_in0</name></connection>
<connection>
<GID>125</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>205,-32,209.5,-32</points>
<connection>
<GID>143</GID>
<name>N_in0</name></connection>
<connection>
<GID>127</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>205,-40,209.5,-40</points>
<connection>
<GID>145</GID>
<name>N_in0</name></connection>
<connection>
<GID>129</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>182,-34,182,-11</points>
<connection>
<GID>135</GID>
<name>OUT_0</name></connection>
<intersection>-34 4</intersection>
<intersection>-15 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>182,-15,199,-15</points>
<connection>
<GID>123</GID>
<name>IN_1</name></connection>
<intersection>182 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>182,-34,199,-34</points>
<connection>
<GID>127</GID>
<name>IN_2</name></connection>
<intersection>182 0</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>258,-86,258,-10</points>
<connection>
<GID>158</GID>
<name>IN_0</name></connection>
<connection>
<GID>151</GID>
<name>OUT_0</name></connection>
<intersection>-86 17</intersection>
<intersection>-76 15</intersection>
<intersection>-66 13</intersection>
<intersection>-46 11</intersection>
<intersection>-36 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>258,-36,284,-36</points>
<connection>
<GID>170</GID>
<name>IN_1</name></connection>
<intersection>258 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>258,-46,284,-46</points>
<connection>
<GID>171</GID>
<name>IN_1</name></connection>
<intersection>258 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>258,-66,284,-66</points>
<connection>
<GID>183</GID>
<name>IN_1</name></connection>
<intersection>258 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>258,-76,284,-76</points>
<connection>
<GID>184</GID>
<name>IN_1</name></connection>
<intersection>258 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>258,-86,284,-86</points>
<connection>
<GID>185</GID>
<name>IN_1</name></connection>
<intersection>258 0</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>266.5,-88,266.5,-10</points>
<connection>
<GID>152</GID>
<name>OUT_0</name></connection>
<intersection>-88 12</intersection>
<intersection>-74 10</intersection>
<intersection>-54 8</intersection>
<intersection>-11 13</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>266.5,-54,284,-54</points>
<connection>
<GID>182</GID>
<name>IN_0</name></connection>
<intersection>266.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>266.5,-74,284,-74</points>
<connection>
<GID>184</GID>
<name>IN_0</name></connection>
<intersection>266.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>266.5,-88,284,-88</points>
<connection>
<GID>185</GID>
<name>IN_2</name></connection>
<intersection>266.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>266.5,-11,266.5,-11</points>
<connection>
<GID>159</GID>
<name>IN_0</name></connection>
<intersection>266.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>290,-17,292.5,-17</points>
<connection>
<GID>168</GID>
<name>OUT</name></connection>
<connection>
<GID>160</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>290,-27,292.5,-27</points>
<connection>
<GID>169</GID>
<name>OUT</name></connection>
<connection>
<GID>161</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>290,-37,292.5,-37</points>
<connection>
<GID>170</GID>
<name>OUT</name></connection>
<connection>
<GID>162</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>290,-47,292.5,-47</points>
<connection>
<GID>171</GID>
<name>OUT</name></connection>
<connection>
<GID>163</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>249.5,-84,249.5,-10</points>
<connection>
<GID>173</GID>
<name>IN_0</name></connection>
<connection>
<GID>172</GID>
<name>OUT_0</name></connection>
<intersection>-84 6</intersection>
<intersection>-44 4</intersection>
<intersection>-24 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>249.5,-24,284,-24</points>
<connection>
<GID>169</GID>
<name>IN_0</name></connection>
<intersection>249.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>249.5,-44,284,-44</points>
<connection>
<GID>171</GID>
<name>IN_0</name></connection>
<intersection>249.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>249.5,-84,284,-84</points>
<connection>
<GID>185</GID>
<name>IN_0</name></connection>
<intersection>249.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>253.5,-78,253.5,-11</points>
<connection>
<GID>173</GID>
<name>OUT_0</name></connection>
<intersection>-78 10</intersection>
<intersection>-64 8</intersection>
<intersection>-58 6</intersection>
<intersection>-34 4</intersection>
<intersection>-14 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>253.5,-14,284,-14</points>
<connection>
<GID>168</GID>
<name>IN_0</name></connection>
<intersection>253.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>253.5,-34,284,-34</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<intersection>253.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>253.5,-58,284,-58</points>
<connection>
<GID>182</GID>
<name>IN_2</name></connection>
<intersection>253.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>253.5,-64,284,-64</points>
<connection>
<GID>183</GID>
<name>IN_0</name></connection>
<intersection>253.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>253.5,-78,284,-78</points>
<connection>
<GID>184</GID>
<name>IN_2</name></connection>
<intersection>253.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>262,-56,262,-11</points>
<connection>
<GID>158</GID>
<name>OUT_0</name></connection>
<intersection>-56 6</intersection>
<intersection>-26 4</intersection>
<intersection>-16 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>262,-16,284,-16</points>
<connection>
<GID>168</GID>
<name>IN_1</name></connection>
<intersection>262 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>262,-26,284,-26</points>
<connection>
<GID>169</GID>
<name>IN_1</name></connection>
<intersection>262 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>262,-56,284,-56</points>
<connection>
<GID>182</GID>
<name>IN_1</name></connection>
<intersection>262 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>270.5,-68,270.5,-11</points>
<connection>
<GID>159</GID>
<name>OUT_0</name></connection>
<intersection>-68 10</intersection>
<intersection>-48 8</intersection>
<intersection>-38 6</intersection>
<intersection>-28 4</intersection>
<intersection>-18 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>270.5,-18,284,-18</points>
<connection>
<GID>168</GID>
<name>IN_2</name></connection>
<intersection>270.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>270.5,-28,284,-28</points>
<connection>
<GID>169</GID>
<name>IN_2</name></connection>
<intersection>270.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>270.5,-38,284,-38</points>
<connection>
<GID>170</GID>
<name>IN_2</name></connection>
<intersection>270.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>270.5,-48,284,-48</points>
<connection>
<GID>171</GID>
<name>IN_2</name></connection>
<intersection>270.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>270.5,-68,284,-68</points>
<connection>
<GID>183</GID>
<name>IN_2</name></connection>
<intersection>270.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274,-90,274,-10</points>
<connection>
<GID>153</GID>
<name>OUT_0</name></connection>
<intersection>-90 13</intersection>
<intersection>-80 14</intersection>
<intersection>-70 11</intersection>
<intersection>-60 9</intersection>
<intersection>-50 7</intersection>
<intersection>-40 5</intersection>
<intersection>-30 3</intersection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>274,-20,284,-20</points>
<connection>
<GID>168</GID>
<name>IN_3</name></connection>
<intersection>274 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>274,-30,284,-30</points>
<connection>
<GID>169</GID>
<name>IN_3</name></connection>
<intersection>274 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>274,-40,284,-40</points>
<connection>
<GID>170</GID>
<name>IN_3</name></connection>
<intersection>274 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>274,-50,284,-50</points>
<connection>
<GID>171</GID>
<name>IN_3</name></connection>
<intersection>274 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>274,-60,284,-60</points>
<connection>
<GID>182</GID>
<name>IN_3</name></connection>
<intersection>274 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>274,-70,284,-70</points>
<connection>
<GID>183</GID>
<name>IN_3</name></connection>
<intersection>274 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>274,-90,284,-90</points>
<connection>
<GID>185</GID>
<name>IN_3</name></connection>
<intersection>274 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>274,-80,284,-80</points>
<connection>
<GID>184</GID>
<name>IN_3</name></connection>
<intersection>274 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>290,-57,292.5,-57</points>
<connection>
<GID>182</GID>
<name>OUT</name></connection>
<connection>
<GID>178</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>290,-67,292.5,-67</points>
<connection>
<GID>183</GID>
<name>OUT</name></connection>
<connection>
<GID>179</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>290,-77,292.5,-77</points>
<connection>
<GID>184</GID>
<name>OUT</name></connection>
<connection>
<GID>180</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>290,-87,292.5,-87</points>
<connection>
<GID>185</GID>
<name>OUT</name></connection>
<connection>
<GID>181</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>362,-43,362,-10</points>
<connection>
<GID>197</GID>
<name>OUT_0</name></connection>
<intersection>-43 4</intersection>
<intersection>-31 3</intersection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>362,-19,368,-19</points>
<connection>
<GID>199</GID>
<name>IN_3</name></connection>
<intersection>362 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>362,-31,368,-31</points>
<connection>
<GID>200</GID>
<name>IN_3</name></connection>
<intersection>362 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>362,-43,368,-43</points>
<connection>
<GID>201</GID>
<name>IN_3</name></connection>
<intersection>362 0</intersection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>357,-29,357,-10</points>
<connection>
<GID>196</GID>
<name>OUT_0</name></connection>
<intersection>-29 3</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>357,-17,368,-17</points>
<connection>
<GID>199</GID>
<name>IN_2</name></connection>
<intersection>357 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>357,-29,368,-29</points>
<connection>
<GID>200</GID>
<name>IN_2</name></connection>
<intersection>357 0</intersection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>352,-41,352,-10</points>
<connection>
<GID>195</GID>
<name>OUT_0</name></connection>
<intersection>-41 2</intersection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>352,-15,368,-15</points>
<connection>
<GID>199</GID>
<name>IN_1</name></connection>
<intersection>352 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>352,-41,368,-41</points>
<connection>
<GID>201</GID>
<name>IN_2</name></connection>
<intersection>352 0</intersection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>347,-13,347,-10</points>
<connection>
<GID>194</GID>
<name>OUT_0</name></connection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>347,-13,368,-13</points>
<connection>
<GID>199</GID>
<name>IN_0</name></connection>
<intersection>347 0</intersection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>337,-25,337,-10</points>
<connection>
<GID>192</GID>
<name>OUT_0</name></connection>
<intersection>-25 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>337,-25,368,-25</points>
<connection>
<GID>200</GID>
<name>IN_0</name></connection>
<intersection>337 0</intersection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>342,-39,342,-10</points>
<connection>
<GID>193</GID>
<name>OUT_0</name></connection>
<intersection>-39 2</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>342,-27,368,-27</points>
<connection>
<GID>200</GID>
<name>IN_1</name></connection>
<intersection>342 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>342,-39,368,-39</points>
<connection>
<GID>201</GID>
<name>IN_1</name></connection>
<intersection>342 0</intersection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>332,-37,332,-10</points>
<connection>
<GID>190</GID>
<name>OUT_0</name></connection>
<intersection>-37 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>332,-37,368,-37</points>
<connection>
<GID>201</GID>
<name>IN_0</name></connection>
<intersection>332 0</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>375,-16,378,-16</points>
<connection>
<GID>203</GID>
<name>N_in0</name></connection>
<connection>
<GID>199</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>375,-28,378,-28</points>
<connection>
<GID>205</GID>
<name>N_in0</name></connection>
<connection>
<GID>200</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>375,-40,378,-40</points>
<connection>
<GID>207</GID>
<name>N_in0</name></connection>
<connection>
<GID>201</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 1>
<page 2>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 2>
<page 3>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 3>
<page 4>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 4>
<page 5>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 5>
<page 6>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 6>
<page 7>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 7>
<page 8>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 9></circuit>