<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-158.955,55.5518,123.188,-83.9061</PageViewport>
<gate>
<ID>41</ID>
<type>AA_AND2</type>
<position>-93,49</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_TOGGLE</type>
<position>-105,51</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>43</ID>
<type>AA_TOGGLE</type>
<position>-105,47.5</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>44</ID>
<type>GA_LED</type>
<position>-87,49</position>
<input>
<ID>N_in0</ID>12 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>45</ID>
<type>AA_LABEL</type>
<position>-122,50</position>
<gparam>LABEL_TEXT AND Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>46</ID>
<type>AA_LABEL</type>
<position>-110,51.5</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>47</ID>
<type>AA_LABEL</type>
<position>-110,47.5</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>AA_LABEL</type>
<position>-78.5,49.5</position>
<gparam>LABEL_TEXT Y = A . B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>49</ID>
<type>AE_OR2</type>
<position>-93,38.5</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_TOGGLE</type>
<position>-105,41</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>51</ID>
<type>AA_TOGGLE</type>
<position>-105,36.5</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>52</ID>
<type>GA_LED</type>
<position>-87,38.5</position>
<input>
<ID>N_in0</ID>15 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>53</ID>
<type>AA_LABEL</type>
<position>-110,41</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>54</ID>
<type>AA_LABEL</type>
<position>-110,37</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>55</ID>
<type>AA_LABEL</type>
<position>-77.5,39</position>
<gparam>LABEL_TEXT Y = A + B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>56</ID>
<type>AI_XOR2</type>
<position>-93,29</position>
<input>
<ID>IN_0</ID>16 </input>
<input>
<ID>IN_1</ID>17 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>57</ID>
<type>AA_TOGGLE</type>
<position>-105,31</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>58</ID>
<type>AA_TOGGLE</type>
<position>-105,27</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>59</ID>
<type>GA_LED</type>
<position>-87,29</position>
<input>
<ID>N_in0</ID>18 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>AA_LABEL</type>
<position>-74.5,29.5</position>
<gparam>LABEL_TEXT Y = A'B + B'A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>61</ID>
<type>AA_LABEL</type>
<position>-122,39.5</position>
<gparam>LABEL_TEXT OR Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>62</ID>
<type>AA_LABEL</type>
<position>-121.5,29</position>
<gparam>LABEL_TEXT XOR Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>64</ID>
<type>AO_XNOR2</type>
<position>-93,19</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>20 </input>
<output>
<ID>OUT</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>66</ID>
<type>AA_TOGGLE</type>
<position>-105,21</position>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>68</ID>
<type>AA_TOGGLE</type>
<position>-105,17</position>
<output>
<ID>OUT_0</ID>20 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>70</ID>
<type>GA_LED</type>
<position>-87,19</position>
<input>
<ID>N_in0</ID>21 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>71</ID>
<type>AA_LABEL</type>
<position>-74,19.5</position>
<gparam>LABEL_TEXT Y = AB + A'B'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>72</ID>
<type>AA_LABEL</type>
<position>-110,21</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>73</ID>
<type>AA_LABEL</type>
<position>-110,17</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>74</ID>
<type>AA_LABEL</type>
<position>-122.5,19.5</position>
<gparam>LABEL_TEXT XNOR Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>76</ID>
<type>BA_NAND2</type>
<position>-93,10</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>23 </input>
<output>
<ID>OUT</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>78</ID>
<type>AA_TOGGLE</type>
<position>-105,12</position>
<output>
<ID>OUT_0</ID>22 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>80</ID>
<type>AA_TOGGLE</type>
<position>-105,8</position>
<output>
<ID>OUT_0</ID>23 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>82</ID>
<type>GA_LED</type>
<position>-87,10</position>
<input>
<ID>N_in0</ID>24 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>83</ID>
<type>AA_LABEL</type>
<position>-76,10.5</position>
<gparam>LABEL_TEXT Y = (A*B)'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>84</ID>
<type>AA_LABEL</type>
<position>-122.5,11</position>
<gparam>LABEL_TEXT Nand Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>85</ID>
<type>AA_LABEL</type>
<position>-110,31</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>86</ID>
<type>AA_LABEL</type>
<position>-110,27</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>87</ID>
<type>AA_LABEL</type>
<position>-110,12</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>88</ID>
<type>AA_LABEL</type>
<position>-110,8</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>90</ID>
<type>BE_NOR2</type>
<position>-93,1</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>92</ID>
<type>AA_TOGGLE</type>
<position>-105,3</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>94</ID>
<type>AA_TOGGLE</type>
<position>-105,-1</position>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>96</ID>
<type>GA_LED</type>
<position>-87,1</position>
<input>
<ID>N_in0</ID>27 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>97</ID>
<type>AA_LABEL</type>
<position>-75.5,1.5</position>
<gparam>LABEL_TEXT Y = (A+B)'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>98</ID>
<type>AA_LABEL</type>
<position>-122,1</position>
<gparam>LABEL_TEXT NOR Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>100</ID>
<type>AA_INVERTER</type>
<position>-93,-7</position>
<input>
<ID>IN_0</ID>28 </input>
<output>
<ID>OUT_0</ID>29 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>102</ID>
<type>AA_TOGGLE</type>
<position>-105,-7</position>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>104</ID>
<type>GA_LED</type>
<position>-87,-7</position>
<input>
<ID>N_in0</ID>29 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>105</ID>
<type>AA_LABEL</type>
<position>-79,-6.5</position>
<gparam>LABEL_TEXT Y = A'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>106</ID>
<type>AA_LABEL</type>
<position>-110,3.5</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>107</ID>
<type>AA_LABEL</type>
<position>-110,-0.5</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>108</ID>
<type>AA_LABEL</type>
<position>-110,-6.5</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>109</ID>
<type>AA_LABEL</type>
<position>-122.5,-6</position>
<gparam>LABEL_TEXT NOT Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-103,51,-96,51</points>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<intersection>-96 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-96,50,-96,51</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<intersection>51 1</intersection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-96.5,47.5,-96.5,48</points>
<intersection>47.5 1</intersection>
<intersection>48 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-103,47.5,-96.5,47.5</points>
<connection>
<GID>43</GID>
<name>OUT_0</name></connection>
<intersection>-96.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-96.5,48,-96,48</points>
<connection>
<GID>41</GID>
<name>IN_1</name></connection>
<intersection>-96.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-90,49,-88,49</points>
<connection>
<GID>41</GID>
<name>OUT</name></connection>
<connection>
<GID>44</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-96,39.5,-96,41</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<intersection>41 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-103,41,-96,41</points>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection>
<intersection>-96 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-96,36.5,-96,37.5</points>
<connection>
<GID>49</GID>
<name>IN_1</name></connection>
<intersection>36.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-103,36.5,-96,36.5</points>
<connection>
<GID>51</GID>
<name>OUT_0</name></connection>
<intersection>-96 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-90,38.5,-88,38.5</points>
<connection>
<GID>49</GID>
<name>OUT</name></connection>
<connection>
<GID>52</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-96,30,-96,31</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>31 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-103,31,-96,31</points>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection>
<intersection>-96 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-96,27,-96,28</points>
<connection>
<GID>56</GID>
<name>IN_1</name></connection>
<intersection>27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-103,27,-96,27</points>
<connection>
<GID>58</GID>
<name>OUT_0</name></connection>
<intersection>-96 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-90,29,-88,29</points>
<connection>
<GID>56</GID>
<name>OUT</name></connection>
<connection>
<GID>59</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-96,20,-96,21</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-103,21,-96,21</points>
<connection>
<GID>66</GID>
<name>OUT_0</name></connection>
<intersection>-96 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-96,17,-96,18</points>
<connection>
<GID>64</GID>
<name>IN_1</name></connection>
<intersection>17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-103,17,-96,17</points>
<connection>
<GID>68</GID>
<name>OUT_0</name></connection>
<intersection>-96 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-90,19,-88,19</points>
<connection>
<GID>64</GID>
<name>OUT</name></connection>
<connection>
<GID>70</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-96,11,-96,12</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-103,12,-96,12</points>
<connection>
<GID>78</GID>
<name>OUT_0</name></connection>
<intersection>-96 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-96,8,-96,9</points>
<connection>
<GID>76</GID>
<name>IN_1</name></connection>
<intersection>8 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-103,8,-96,8</points>
<connection>
<GID>80</GID>
<name>OUT_0</name></connection>
<intersection>-96 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-90,10,-88,10</points>
<connection>
<GID>82</GID>
<name>N_in0</name></connection>
<connection>
<GID>76</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-96,2,-96,3</points>
<connection>
<GID>90</GID>
<name>IN_0</name></connection>
<intersection>3 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-103,3,-96,3</points>
<connection>
<GID>92</GID>
<name>OUT_0</name></connection>
<intersection>-96 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-96,-1,-96,0</points>
<connection>
<GID>90</GID>
<name>IN_1</name></connection>
<intersection>-1 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-103,-1,-96,-1</points>
<connection>
<GID>94</GID>
<name>OUT_0</name></connection>
<intersection>-96 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-90,1,-88,1</points>
<connection>
<GID>90</GID>
<name>OUT</name></connection>
<connection>
<GID>96</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-103,-7,-96,-7</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<connection>
<GID>102</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-90,-7,-88,-7</points>
<connection>
<GID>100</GID>
<name>OUT_0</name></connection>
<connection>
<GID>104</GID>
<name>N_in0</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>606.697,-22.0445,675.624,-56.1142</PageViewport>
<gate>
<ID>193</ID>
<type>AA_LABEL</type>
<position>391.5,-64.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1</ID>
<type>AA_LABEL</type>
<position>104.5,-36.5</position>
<gparam>LABEL_TEXT Y = (A*B)</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>194</ID>
<type>AA_TOGGLE</type>
<position>375,-30.5</position>
<output>
<ID>OUT_0</ID>94 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>195</ID>
<type>AA_LABEL</type>
<position>528,-13</position>
<gparam>LABEL_TEXT Half Adder NAND Implementation</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2</ID>
<type>AA_LABEL</type>
<position>109,-48.5</position>
<gparam>LABEL_TEXT Y = (A+B)</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3</ID>
<type>AA_LABEL</type>
<position>47,-48.5</position>
<gparam>LABEL_TEXT NAND as a OR Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>196</ID>
<type>AA_AND2</type>
<position>426,-37.5</position>
<input>
<ID>IN_0</ID>93 </input>
<input>
<ID>IN_1</ID>94 </input>
<output>
<ID>OUT</ID>90 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>BA_NAND2</type>
<position>82.5,-62.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_TOGGLE</type>
<position>73.5,-62.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>198</ID>
<type>AA_AND2</type>
<position>426,-43.5</position>
<input>
<ID>IN_0</ID>92 </input>
<input>
<ID>IN_1</ID>95 </input>
<output>
<ID>OUT</ID>91 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>199</ID>
<type>AA_TOGGLE</type>
<position>499.5,-30.5</position>
<output>
<ID>OUT_0</ID>75 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_LABEL</type>
<position>69,-62</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>7</ID>
<type>BA_NAND2</type>
<position>82.5,-70.5</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>200</ID>
<type>AE_OR2</type>
<position>438,-41</position>
<input>
<ID>IN_0</ID>90 </input>
<input>
<ID>IN_1</ID>91 </input>
<output>
<ID>OUT</ID>97 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>74,-70.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_LABEL</type>
<position>69,-70.5</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>202</ID>
<type>AE_SMALL_INVERTER</type>
<position>366.5,-36.5</position>
<input>
<ID>IN_0</ID>92 </input>
<output>
<ID>OUT_0</ID>93 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>203</ID>
<type>AA_TOGGLE</type>
<position>509.5,-30.5</position>
<output>
<ID>OUT_0</ID>76 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>10</ID>
<type>BA_NAND2</type>
<position>93,-66.5</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>204</ID>
<type>AE_SMALL_INVERTER</type>
<position>377,-44.5</position>
<input>
<ID>IN_0</ID>94 </input>
<output>
<ID>OUT_0</ID>95 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>12</ID>
<type>BA_NAND2</type>
<position>101,-66.5</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>205</ID>
<type>AA_AND2</type>
<position>426,-50.5</position>
<input>
<ID>IN_0</ID>92 </input>
<input>
<ID>IN_1</ID>94 </input>
<output>
<ID>OUT</ID>96 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>13</ID>
<type>AI_XOR2</type>
<position>409,-73</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>14</ID>
<type>GA_LED</type>
<position>106,-66.5</position>
<input>
<ID>N_in0</ID>6 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>207</ID>
<type>GA_LED</type>
<position>433,-50.5</position>
<input>
<ID>N_in0</ID>96 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>208</ID>
<type>BA_NAND2</type>
<position>526,-39.5</position>
<input>
<ID>IN_0</ID>60 </input>
<input>
<ID>IN_1</ID>76 </input>
<output>
<ID>OUT</ID>80 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>15</ID>
<type>AA_LABEL</type>
<position>117.5,-66</position>
<gparam>LABEL_TEXT Y = (A+B)'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>AA_LABEL</type>
<position>47,-66</position>
<gparam>LABEL_TEXT NAND as a NOR Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>209</ID>
<type>GA_LED</type>
<position>443.5,-41</position>
<input>
<ID>N_in0</ID>97 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>17</ID>
<type>BA_NAND2</type>
<position>95,-81</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>33 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>BA_NAND2</type>
<position>95,-87</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>211</ID>
<type>AA_LABEL</type>
<position>447.5,-40.5</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>212</ID>
<type>BA_NAND2</type>
<position>526,-47.5</position>
<input>
<ID>IN_0</ID>75 </input>
<input>
<ID>IN_1</ID>78 </input>
<output>
<ID>OUT</ID>98 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>19</ID>
<type>BA_NAND2</type>
<position>84,-84</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_TOGGLE</type>
<position>74,-80</position>
<output>
<ID>OUT_0</ID>31 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>213</ID>
<type>AA_LABEL</type>
<position>441,-50</position>
<gparam>LABEL_TEXT C = AB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>21</ID>
<type>AA_TOGGLE</type>
<position>74,-88</position>
<output>
<ID>OUT_0</ID>32 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>22</ID>
<type>BA_NAND2</type>
<position>104,-84</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>35 </input>
<output>
<ID>OUT</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>215</ID>
<type>AA_LABEL</type>
<position>364.5,-25.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>216</ID>
<type>AE_SMALL_INVERTER</type>
<position>501.5,-38.5</position>
<input>
<ID>IN_0</ID>75 </input>
<output>
<ID>OUT_0</ID>60 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>24</ID>
<type>GA_LED</type>
<position>110,-84</position>
<input>
<ID>N_in0</ID>36 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>217</ID>
<type>AA_LABEL</type>
<position>375,-25.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>25</ID>
<type>AA_AND2</type>
<position>409.5,-80.5</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>56 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>219</ID>
<type>AE_SMALL_INVERTER</type>
<position>511.5,-48.5</position>
<input>
<ID>IN_0</ID>76 </input>
<output>
<ID>OUT_0</ID>78 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_LABEL</type>
<position>123.5,-83.5</position>
<gparam>LABEL_TEXT Y = A'B + B'A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>27</ID>
<type>AA_LABEL</type>
<position>47.5,-84</position>
<gparam>LABEL_TEXT NAND as a XOR Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>221</ID>
<type>BA_NAND2</type>
<position>534.5,-43.5</position>
<input>
<ID>IN_0</ID>80 </input>
<input>
<ID>IN_1</ID>98 </input>
<output>
<ID>OUT</ID>99 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_LABEL</type>
<position>68.5,-79.5</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>29</ID>
<type>AA_LABEL</type>
<position>69,-88</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>223</ID>
<type>GA_LED</type>
<position>540.5,-43.5</position>
<input>
<ID>N_in0</ID>99 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>BA_NAND2</type>
<position>95,-97.5</position>
<input>
<ID>IN_0</ID>37 </input>
<input>
<ID>IN_1</ID>46 </input>
<output>
<ID>OUT</ID>47 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>31</ID>
<type>BA_NAND2</type>
<position>95,-103.5</position>
<input>
<ID>IN_0</ID>46 </input>
<input>
<ID>IN_1</ID>45 </input>
<output>
<ID>OUT</ID>48 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>225</ID>
<type>AA_LABEL</type>
<position>499.5,-25.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>BA_NAND2</type>
<position>84,-100.5</position>
<input>
<ID>IN_0</ID>37 </input>
<input>
<ID>IN_1</ID>45 </input>
<output>
<ID>OUT</ID>46 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>33</ID>
<type>AA_TOGGLE</type>
<position>74,-96.5</position>
<output>
<ID>OUT_0</ID>37 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>227</ID>
<type>AA_LABEL</type>
<position>509.5,-25.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>AA_TOGGLE</type>
<position>74,-104.5</position>
<output>
<ID>OUT_0</ID>45 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>35</ID>
<type>BA_NAND2</type>
<position>104,-100.5</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>48 </input>
<output>
<ID>OUT</ID>49 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>229</ID>
<type>AA_LABEL</type>
<position>546,-43</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>AA_LABEL</type>
<position>68.5,-96</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>230</ID>
<type>BA_NAND2</type>
<position>526,-54.5</position>
<input>
<ID>IN_0</ID>75 </input>
<input>
<ID>IN_1</ID>76 </input>
<output>
<ID>OUT</ID>101 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>37</ID>
<type>AA_LABEL</type>
<position>69,-104.5</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>231</ID>
<type>GA_LED</type>
<position>540,-54.5</position>
<input>
<ID>N_in0</ID>102 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>BA_NAND2</type>
<position>112.5,-100.5</position>
<input>
<ID>IN_0</ID>49 </input>
<input>
<ID>IN_1</ID>49 </input>
<output>
<ID>OUT</ID>53 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>232</ID>
<type>BA_NAND2</type>
<position>534,-54.5</position>
<input>
<ID>IN_0</ID>101 </input>
<input>
<ID>IN_1</ID>101 </input>
<output>
<ID>OUT</ID>102 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>39</ID>
<type>GA_LED</type>
<position>119,-100.5</position>
<input>
<ID>N_in0</ID>53 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>233</ID>
<type>AA_LABEL</type>
<position>545.5,-54</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>AA_LABEL</type>
<position>134,-100</position>
<gparam>LABEL_TEXT Y = AB + A'B'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>234</ID>
<type>AA_LABEL</type>
<position>653,-13</position>
<gparam>LABEL_TEXT Half Adder NOR Implementation</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>236</ID>
<type>AA_TOGGLE</type>
<position>616.5,-24.5</position>
<output>
<ID>OUT_0</ID>103 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>238</ID>
<type>AA_TOGGLE</type>
<position>628.5,-24.5</position>
<output>
<ID>OUT_0</ID>104 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>240</ID>
<type>BE_NOR2</type>
<position>650.5,-31.5</position>
<input>
<ID>IN_0</ID>103 </input>
<input>
<ID>IN_1</ID>105 </input>
<output>
<ID>OUT</ID>107 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>242</ID>
<type>BE_NOR2</type>
<position>650.5,-38.5</position>
<input>
<ID>IN_0</ID>106 </input>
<input>
<ID>IN_1</ID>104 </input>
<output>
<ID>OUT</ID>108 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>244</ID>
<type>AE_SMALL_INVERTER</type>
<position>630.5,-32.5</position>
<input>
<ID>IN_0</ID>104 </input>
<output>
<ID>OUT_0</ID>105 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>246</ID>
<type>AE_SMALL_INVERTER</type>
<position>618.5,-37.5</position>
<input>
<ID>IN_0</ID>103 </input>
<output>
<ID>OUT_0</ID>106 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>248</ID>
<type>BE_NOR2</type>
<position>660.5,-35</position>
<input>
<ID>IN_0</ID>107 </input>
<input>
<ID>IN_1</ID>108 </input>
<output>
<ID>OUT</ID>109 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>250</ID>
<type>BE_NOR2</type>
<position>669,-35</position>
<input>
<ID>IN_0</ID>109 </input>
<input>
<ID>IN_1</ID>109 </input>
<output>
<ID>OUT</ID>110 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>252</ID>
<type>GA_LED</type>
<position>675,-35</position>
<input>
<ID>N_in0</ID>110 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>254</ID>
<type>BE_NOR2</type>
<position>651,-45</position>
<input>
<ID>IN_0</ID>105 </input>
<input>
<ID>IN_1</ID>106 </input>
<output>
<ID>OUT</ID>111 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>256</ID>
<type>BE_NOR2</type>
<position>659.5,-45</position>
<input>
<ID>IN_0</ID>111 </input>
<input>
<ID>IN_1</ID>111 </input>
<output>
<ID>OUT</ID>112 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>63</ID>
<type>AA_LABEL</type>
<position>46.5,-100</position>
<gparam>LABEL_TEXT NAND as a XNOR Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>258</ID>
<type>GA_LED</type>
<position>666,-45</position>
<input>
<ID>N_in0</ID>112 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>65</ID>
<type>AA_LABEL</type>
<position>272,-13.5</position>
<gparam>LABEL_TEXT NOR as a Universal Gate</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>69</ID>
<type>BE_NOR2</type>
<position>272.5,-25.5</position>
<input>
<ID>IN_0</ID>54 </input>
<input>
<ID>IN_1</ID>54 </input>
<output>
<ID>OUT</ID>55 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>75</ID>
<type>AA_TOGGLE</type>
<position>384.5,-68.5</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>77</ID>
<type>AA_TOGGLE</type>
<position>265.5,-25.5</position>
<output>
<ID>OUT_0</ID>54 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>81</ID>
<type>GA_LED</type>
<position>278,-25.5</position>
<input>
<ID>N_in0</ID>55 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>89</ID>
<type>AA_LABEL</type>
<position>262.5,-25</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>91</ID>
<type>AA_LABEL</type>
<position>281,-25</position>
<gparam>LABEL_TEXT A'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>93</ID>
<type>BE_NOR2</type>
<position>272.5,-34.5</position>
<input>
<ID>IN_0</ID>58 </input>
<input>
<ID>IN_1</ID>59 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>95</ID>
<type>BE_NOR2</type>
<position>279.5,-34.5</position>
<input>
<ID>IN_0</ID>57 </input>
<input>
<ID>IN_1</ID>57 </input>
<output>
<ID>OUT</ID>61 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>99</ID>
<type>AA_TOGGLE</type>
<position>265.5,-33</position>
<output>
<ID>OUT_0</ID>58 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>101</ID>
<type>AA_TOGGLE</type>
<position>265.5,-36</position>
<output>
<ID>OUT_0</ID>59 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>103</ID>
<type>AA_TOGGLE</type>
<position>391.5,-68.5</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>110</ID>
<type>AA_LABEL</type>
<position>263,-32.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>111</ID>
<type>AA_LABEL</type>
<position>263,-35.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>113</ID>
<type>AA_LABEL</type>
<position>419,-72.5</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>115</ID>
<type>GA_LED</type>
<position>284.5,-34.5</position>
<input>
<ID>N_in0</ID>61 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>116</ID>
<type>AA_LABEL</type>
<position>288.5,-34</position>
<gparam>LABEL_TEXT A + B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>117</ID>
<type>AA_LABEL</type>
<position>71.5,-13.5</position>
<gparam>LABEL_TEXT NAND as a Universal Gate</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>118</ID>
<type>BE_NOR2</type>
<position>270.5,-42.5</position>
<input>
<ID>IN_0</ID>64 </input>
<input>
<ID>IN_1</ID>64 </input>
<output>
<ID>OUT</ID>62 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>119</ID>
<type>BE_NOR2</type>
<position>270.5,-49.5</position>
<input>
<ID>IN_0</ID>65 </input>
<input>
<ID>IN_1</ID>65 </input>
<output>
<ID>OUT</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>120</ID>
<type>BE_NOR2</type>
<position>278.5,-46</position>
<input>
<ID>IN_0</ID>62 </input>
<input>
<ID>IN_1</ID>63 </input>
<output>
<ID>OUT</ID>66 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>121</ID>
<type>AA_TOGGLE</type>
<position>264,-42.5</position>
<output>
<ID>OUT_0</ID>64 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>122</ID>
<type>AA_TOGGLE</type>
<position>264,-49.5</position>
<output>
<ID>OUT_0</ID>65 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>123</ID>
<type>AA_TOGGLE</type>
<position>76.5,-28</position>
<output>
<ID>OUT_0</ID>38 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>124</ID>
<type>GA_LED</type>
<position>415,-73</position>
<input>
<ID>N_in0</ID>30 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>125</ID>
<type>GA_LED</type>
<position>91.5,-28</position>
<input>
<ID>N_in0</ID>39 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>126</ID>
<type>AA_LABEL</type>
<position>71,-27.5</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>127</ID>
<type>GA_LED</type>
<position>283.5,-46</position>
<input>
<ID>N_in0</ID>66 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>128</ID>
<type>AA_LABEL</type>
<position>288.5,-45.5</position>
<gparam>LABEL_TEXT A . B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>129</ID>
<type>BA_NAND2</type>
<position>84.5,-28</position>
<input>
<ID>IN_0</ID>38 </input>
<input>
<ID>IN_1</ID>38 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>130</ID>
<type>AA_LABEL</type>
<position>101,-27.5</position>
<gparam>LABEL_TEXT Y = A'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>131</ID>
<type>AA_LABEL</type>
<position>48,-27</position>
<gparam>LABEL_TEXT NAND as a NOT Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>132</ID>
<type>BA_NAND2</type>
<position>82,-37</position>
<input>
<ID>IN_0</ID>40 </input>
<input>
<ID>IN_1</ID>41 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>133</ID>
<type>AA_TOGGLE</type>
<position>74,-35</position>
<output>
<ID>OUT_0</ID>40 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>134</ID>
<type>AA_TOGGLE</type>
<position>74,-39</position>
<output>
<ID>OUT_0</ID>41 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>135</ID>
<type>AA_LABEL</type>
<position>69,-34.5</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>136</ID>
<type>AA_LABEL</type>
<position>69,-38.5</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>137</ID>
<type>AA_LABEL</type>
<position>261.5,-42</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>138</ID>
<type>BA_NAND2</type>
<position>89.5,-37</position>
<input>
<ID>IN_0</ID>42 </input>
<input>
<ID>IN_1</ID>42 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>139</ID>
<type>AA_LABEL</type>
<position>261.5,-49</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>140</ID>
<type>GA_LED</type>
<position>94.5,-37</position>
<input>
<ID>N_in0</ID>43 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>141</ID>
<type>AA_LABEL</type>
<position>48,-36.5</position>
<gparam>LABEL_TEXT NAND as a AND Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>142</ID>
<type>BA_NAND2</type>
<position>82.5,-45</position>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_1</ID>44 </input>
<output>
<ID>OUT</ID>50 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>143</ID>
<type>AA_TOGGLE</type>
<position>74,-45</position>
<output>
<ID>OUT_0</ID>44 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>144</ID>
<type>BE_NOR2</type>
<position>270.5,-57</position>
<input>
<ID>IN_0</ID>69 </input>
<input>
<ID>IN_1</ID>69 </input>
<output>
<ID>OUT</ID>67 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>145</ID>
<type>AA_LABEL</type>
<position>69,-44.5</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>146</ID>
<type>BE_NOR2</type>
<position>270.5,-64</position>
<input>
<ID>IN_0</ID>70 </input>
<input>
<ID>IN_1</ID>70 </input>
<output>
<ID>OUT</ID>68 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>147</ID>
<type>BA_NAND2</type>
<position>82.5,-53</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>8 </input>
<output>
<ID>OUT</ID>51 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>148</ID>
<type>AA_TOGGLE</type>
<position>74,-53</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>149</ID>
<type>BE_NOR2</type>
<position>278.5,-60.5</position>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>68 </input>
<output>
<ID>OUT</ID>72 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>150</ID>
<type>AA_TOGGLE</type>
<position>264,-57</position>
<output>
<ID>OUT_0</ID>69 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>151</ID>
<type>AA_LABEL</type>
<position>69,-53</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>152</ID>
<type>BA_NAND2</type>
<position>93,-49</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>51 </input>
<output>
<ID>OUT</ID>52 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>153</ID>
<type>AA_TOGGLE</type>
<position>264,-64</position>
<output>
<ID>OUT_0</ID>70 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>154</ID>
<type>GA_LED</type>
<position>98,-49</position>
<input>
<ID>N_in0</ID>52 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>155</ID>
<type>AA_LABEL</type>
<position>261.5,-56.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>156</ID>
<type>AA_LABEL</type>
<position>261.5,-63.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>157</ID>
<type>BE_NOR2</type>
<position>286,-60.5</position>
<input>
<ID>IN_0</ID>72 </input>
<input>
<ID>IN_1</ID>72 </input>
<output>
<ID>OUT</ID>71 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>158</ID>
<type>GA_LED</type>
<position>291,-60.5</position>
<input>
<ID>N_in0</ID>71 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>159</ID>
<type>AA_LABEL</type>
<position>296,-60</position>
<gparam>LABEL_TEXT (A + B)'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>160</ID>
<type>BE_NOR2</type>
<position>281.5,-74</position>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>79 </input>
<output>
<ID>OUT</ID>73 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>161</ID>
<type>BE_NOR2</type>
<position>281.5,-81</position>
<input>
<ID>IN_0</ID>79 </input>
<input>
<ID>IN_1</ID>82 </input>
<output>
<ID>OUT</ID>74 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>162</ID>
<type>BE_NOR2</type>
<position>289.5,-77.5</position>
<input>
<ID>IN_0</ID>73 </input>
<input>
<ID>IN_1</ID>74 </input>
<output>
<ID>OUT</ID>77 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>163</ID>
<type>BE_NOR2</type>
<position>297,-77.5</position>
<input>
<ID>IN_0</ID>77 </input>
<input>
<ID>IN_1</ID>77 </input>
<output>
<ID>OUT</ID>83 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>164</ID>
<type>BE_NOR2</type>
<position>272.5,-77.5</position>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>82 </input>
<output>
<ID>OUT</ID>79 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>166</ID>
<type>AA_TOGGLE</type>
<position>263.5,-73</position>
<output>
<ID>OUT_0</ID>81 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>167</ID>
<type>AA_TOGGLE</type>
<position>263.5,-82</position>
<output>
<ID>OUT_0</ID>82 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>168</ID>
<type>GA_LED</type>
<position>415,-80.5</position>
<input>
<ID>N_in0</ID>56 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>169</ID>
<type>GA_LED</type>
<position>302.5,-77.5</position>
<input>
<ID>N_in0</ID>83 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>170</ID>
<type>AA_LABEL</type>
<position>308.5,-77</position>
<gparam>LABEL_TEXT A'B + AB'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>171</ID>
<type>AA_LABEL</type>
<position>261,-82</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>172</ID>
<type>AA_LABEL</type>
<position>261,-73</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>173</ID>
<type>BE_NOR2</type>
<position>281.5,-90.5</position>
<input>
<ID>IN_0</ID>87 </input>
<input>
<ID>IN_1</ID>86 </input>
<output>
<ID>OUT</ID>84 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>174</ID>
<type>BE_NOR2</type>
<position>281.5,-97.5</position>
<input>
<ID>IN_0</ID>86 </input>
<input>
<ID>IN_1</ID>88 </input>
<output>
<ID>OUT</ID>85 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>175</ID>
<type>BE_NOR2</type>
<position>289.5,-94</position>
<input>
<ID>IN_0</ID>84 </input>
<input>
<ID>IN_1</ID>85 </input>
<output>
<ID>OUT</ID>89 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>176</ID>
<type>BE_NOR2</type>
<position>272.5,-94</position>
<input>
<ID>IN_0</ID>87 </input>
<input>
<ID>IN_1</ID>88 </input>
<output>
<ID>OUT</ID>86 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>177</ID>
<type>AA_TOGGLE</type>
<position>263.5,-89.5</position>
<output>
<ID>OUT_0</ID>87 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>178</ID>
<type>AA_TOGGLE</type>
<position>263.5,-98.5</position>
<output>
<ID>OUT_0</ID>88 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>179</ID>
<type>AA_LABEL</type>
<position>261,-98.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>180</ID>
<type>AA_LABEL</type>
<position>261,-89.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>181</ID>
<type>AA_LABEL</type>
<position>419,-80</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>182</ID>
<type>GA_LED</type>
<position>295,-94</position>
<input>
<ID>N_in0</ID>89 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>183</ID>
<type>AA_LABEL</type>
<position>301,-93.5</position>
<gparam>LABEL_TEXT AB + A'B'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>184</ID>
<type>AA_LABEL</type>
<position>243.5,-24.5</position>
<gparam>LABEL_TEXT NOR as a NOT Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>185</ID>
<type>AA_LABEL</type>
<position>243,-33.5</position>
<gparam>LABEL_TEXT NOR as a OR Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>186</ID>
<type>AA_LABEL</type>
<position>243,-45</position>
<gparam>LABEL_TEXT NOR as a AND Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>187</ID>
<type>AA_LABEL</type>
<position>243,-60.5</position>
<gparam>LABEL_TEXT NOR as a NAND Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>188</ID>
<type>AA_LABEL</type>
<position>243,-76.5</position>
<gparam>LABEL_TEXT NOR as a XOR Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>189</ID>
<type>AA_LABEL</type>
<position>244,-93.5</position>
<gparam>LABEL_TEXT NOR as a XNOR Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>190</ID>
<type>AA_LABEL</type>
<position>413.5,-13.5</position>
<gparam>LABEL_TEXT Half Adder</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>191</ID>
<type>AA_LABEL</type>
<position>384.5,-64.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>192</ID>
<type>AA_TOGGLE</type>
<position>364.5,-30.5</position>
<output>
<ID>OUT_0</ID>92 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78,-63.5,78,-61.5</points>
<intersection>-63.5 4</intersection>
<intersection>-62.5 3</intersection>
<intersection>-61.5 5</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75.5,-62.5,78,-62.5</points>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection>
<intersection>78 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>78,-63.5,79.5,-63.5</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>78 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>78,-61.5,79.5,-61.5</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>78 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,-70.5,78,-70.5</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>78 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>78,-71.5,78,-69.5</points>
<intersection>-71.5 10</intersection>
<intersection>-70.5 1</intersection>
<intersection>-69.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>78,-69.5,79.5,-69.5</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>78 8</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>78,-71.5,79.5,-71.5</points>
<connection>
<GID>7</GID>
<name>IN_1</name></connection>
<intersection>78 8</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87.5,-65.5,87.5,-62.5</points>
<intersection>-65.5 2</intersection>
<intersection>-62.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85.5,-62.5,87.5,-62.5</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<intersection>87.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>87.5,-65.5,90,-65.5</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>87.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87.5,-70.5,87.5,-67.5</points>
<intersection>-70.5 1</intersection>
<intersection>-67.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85.5,-70.5,87.5,-70.5</points>
<connection>
<GID>7</GID>
<name>OUT</name></connection>
<intersection>87.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>87.5,-67.5,90,-67.5</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<intersection>87.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97,-67.5,97,-65.5</points>
<intersection>-67.5 3</intersection>
<intersection>-66.5 1</intersection>
<intersection>-65.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>96,-66.5,97,-66.5</points>
<connection>
<GID>10</GID>
<name>OUT</name></connection>
<intersection>97 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97,-65.5,98,-65.5</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>97 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>97,-67.5,98,-67.5</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<intersection>97 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104,-66.5,105,-66.5</points>
<connection>
<GID>12</GID>
<name>OUT</name></connection>
<connection>
<GID>14</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>384.5,-79.5,384.5,-70.5</points>
<connection>
<GID>75</GID>
<name>OUT_0</name></connection>
<intersection>-79.5 3</intersection>
<intersection>-72 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>384.5,-72,406,-72</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<intersection>384.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>384.5,-79.5,406.5,-79.5</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>384.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,-53,78,-53</points>
<connection>
<GID>148</GID>
<name>OUT_0</name></connection>
<intersection>78 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>78,-54,78,-52</points>
<intersection>-54 4</intersection>
<intersection>-53 1</intersection>
<intersection>-52 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>78,-54,79.5,-54</points>
<connection>
<GID>147</GID>
<name>IN_1</name></connection>
<intersection>78 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>78,-52,79.5,-52</points>
<connection>
<GID>147</GID>
<name>IN_0</name></connection>
<intersection>78 3</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>391.5,-81.5,391.5,-70.5</points>
<connection>
<GID>103</GID>
<name>OUT_0</name></connection>
<intersection>-81.5 3</intersection>
<intersection>-74 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>391.5,-74,406,-74</points>
<connection>
<GID>13</GID>
<name>IN_1</name></connection>
<intersection>391.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>391.5,-81.5,406.5,-81.5</points>
<connection>
<GID>25</GID>
<name>IN_1</name></connection>
<intersection>391.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>412,-73,414,-73</points>
<connection>
<GID>13</GID>
<name>OUT</name></connection>
<connection>
<GID>124</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,-80,92,-80</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>78.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>78.5,-83,78.5,-80</points>
<intersection>-83 5</intersection>
<intersection>-80 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>78.5,-83,81,-83</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>78.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,-88,92,-88</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<connection>
<GID>21</GID>
<name>OUT_0</name></connection>
<intersection>78.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>78.5,-88,78.5,-85</points>
<intersection>-88 1</intersection>
<intersection>-85 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>78.5,-85,81,-85</points>
<connection>
<GID>19</GID>
<name>IN_1</name></connection>
<intersection>78.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-86,89.5,-82</points>
<intersection>-86 3</intersection>
<intersection>-84 1</intersection>
<intersection>-82 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>87,-84,89.5,-84</points>
<connection>
<GID>19</GID>
<name>OUT</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>89.5,-82,92,-82</points>
<connection>
<GID>17</GID>
<name>IN_1</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>89.5,-86,92,-86</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99.5,-83,99.5,-81</points>
<intersection>-83 1</intersection>
<intersection>-81 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99.5,-83,101,-83</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>99.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>98,-81,99.5,-81</points>
<connection>
<GID>17</GID>
<name>OUT</name></connection>
<intersection>99.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99.5,-87,99.5,-85</points>
<intersection>-87 2</intersection>
<intersection>-85 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99.5,-85,101,-85</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>99.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>98,-87,99.5,-87</points>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<intersection>99.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>107,-84,109,-84</points>
<connection>
<GID>22</GID>
<name>OUT</name></connection>
<connection>
<GID>24</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,-96.5,92,-96.5</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<connection>
<GID>33</GID>
<name>OUT_0</name></connection>
<intersection>78.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>78.5,-99.5,78.5,-96.5</points>
<intersection>-99.5 5</intersection>
<intersection>-96.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>78.5,-99.5,81,-99.5</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>78.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-29,80,-27</points>
<intersection>-29 3</intersection>
<intersection>-28 1</intersection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>78.5,-28,80,-28</points>
<connection>
<GID>123</GID>
<name>OUT_0</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>80,-27,81.5,-27</points>
<connection>
<GID>129</GID>
<name>IN_0</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>80,-29,81.5,-29</points>
<connection>
<GID>129</GID>
<name>IN_1</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>87.5,-28,90.5,-28</points>
<connection>
<GID>125</GID>
<name>N_in0</name></connection>
<connection>
<GID>129</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79,-36,79,-35</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76,-35,79,-35</points>
<connection>
<GID>133</GID>
<name>OUT_0</name></connection>
<intersection>79 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79,-39,79,-38</points>
<connection>
<GID>132</GID>
<name>IN_1</name></connection>
<intersection>-39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76,-39,79,-39</points>
<connection>
<GID>134</GID>
<name>OUT_0</name></connection>
<intersection>79 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85.5,-38,85.5,-36</points>
<intersection>-38 3</intersection>
<intersection>-37 2</intersection>
<intersection>-36 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85.5,-36,86.5,-36</points>
<connection>
<GID>138</GID>
<name>IN_0</name></connection>
<intersection>85.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>85,-37,85.5,-37</points>
<connection>
<GID>132</GID>
<name>OUT</name></connection>
<intersection>85.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>85.5,-38,86.5,-38</points>
<connection>
<GID>138</GID>
<name>IN_1</name></connection>
<intersection>85.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>92.5,-37,93.5,-37</points>
<connection>
<GID>138</GID>
<name>OUT</name></connection>
<connection>
<GID>140</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78,-46,78,-44</points>
<intersection>-46 4</intersection>
<intersection>-45 3</intersection>
<intersection>-44 5</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>76,-45,78,-45</points>
<connection>
<GID>143</GID>
<name>OUT_0</name></connection>
<intersection>78 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>78,-46,79.5,-46</points>
<connection>
<GID>142</GID>
<name>IN_1</name></connection>
<intersection>78 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>78,-44,79.5,-44</points>
<connection>
<GID>142</GID>
<name>IN_0</name></connection>
<intersection>78 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,-104.5,92,-104.5</points>
<connection>
<GID>31</GID>
<name>IN_1</name></connection>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection>
<intersection>78.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>78.5,-104.5,78.5,-101.5</points>
<intersection>-104.5 1</intersection>
<intersection>-101.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>78.5,-101.5,81,-101.5</points>
<connection>
<GID>32</GID>
<name>IN_1</name></connection>
<intersection>78.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-102.5,89.5,-98.5</points>
<intersection>-102.5 3</intersection>
<intersection>-100.5 1</intersection>
<intersection>-98.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>87,-100.5,89.5,-100.5</points>
<connection>
<GID>32</GID>
<name>OUT</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>89.5,-98.5,92,-98.5</points>
<connection>
<GID>30</GID>
<name>IN_1</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>89.5,-102.5,92,-102.5</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99.5,-99.5,99.5,-97.5</points>
<intersection>-99.5 1</intersection>
<intersection>-97.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99.5,-99.5,101,-99.5</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<intersection>99.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>98,-97.5,99.5,-97.5</points>
<connection>
<GID>30</GID>
<name>OUT</name></connection>
<intersection>99.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99.5,-103.5,99.5,-101.5</points>
<intersection>-103.5 2</intersection>
<intersection>-101.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99.5,-101.5,101,-101.5</points>
<connection>
<GID>35</GID>
<name>IN_1</name></connection>
<intersection>99.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>98,-103.5,99.5,-103.5</points>
<connection>
<GID>31</GID>
<name>OUT</name></connection>
<intersection>99.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,-101.5,108,-99.5</points>
<intersection>-101.5 3</intersection>
<intersection>-100.5 2</intersection>
<intersection>-99.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108,-99.5,109.5,-99.5</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>108 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>107,-100.5,108,-100.5</points>
<connection>
<GID>35</GID>
<name>OUT</name></connection>
<intersection>108 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>108,-101.5,109.5,-101.5</points>
<connection>
<GID>38</GID>
<name>IN_1</name></connection>
<intersection>108 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87.5,-48,87.5,-45</points>
<intersection>-48 2</intersection>
<intersection>-45 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85.5,-45,87.5,-45</points>
<connection>
<GID>142</GID>
<name>OUT</name></connection>
<intersection>87.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>87.5,-48,90,-48</points>
<connection>
<GID>152</GID>
<name>IN_0</name></connection>
<intersection>87.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87.5,-53,87.5,-50</points>
<intersection>-53 1</intersection>
<intersection>-50 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85.5,-53,87.5,-53</points>
<connection>
<GID>147</GID>
<name>OUT</name></connection>
<intersection>87.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>87.5,-50,90,-50</points>
<connection>
<GID>152</GID>
<name>IN_1</name></connection>
<intersection>87.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>96,-49,97,-49</points>
<connection>
<GID>152</GID>
<name>OUT</name></connection>
<connection>
<GID>154</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>115.5,-100.5,118,-100.5</points>
<connection>
<GID>38</GID>
<name>OUT</name></connection>
<connection>
<GID>39</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>268.5,-26.5,268.5,-24.5</points>
<intersection>-26.5 3</intersection>
<intersection>-25.5 1</intersection>
<intersection>-24.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>267.5,-25.5,268.5,-25.5</points>
<connection>
<GID>77</GID>
<name>OUT_0</name></connection>
<intersection>268.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>268.5,-24.5,269.5,-24.5</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<intersection>268.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>268.5,-26.5,269.5,-26.5</points>
<connection>
<GID>69</GID>
<name>IN_1</name></connection>
<intersection>268.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>275.5,-25.5,277,-25.5</points>
<connection>
<GID>69</GID>
<name>OUT</name></connection>
<connection>
<GID>81</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>412.5,-80.5,414,-80.5</points>
<connection>
<GID>25</GID>
<name>OUT</name></connection>
<connection>
<GID>168</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>275.5,-35.5,275.5,-33.5</points>
<intersection>-35.5 3</intersection>
<intersection>-33.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>275.5,-33.5,276.5,-33.5</points>
<connection>
<GID>95</GID>
<name>IN_0</name></connection>
<intersection>275.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>275.5,-35.5,276.5,-35.5</points>
<connection>
<GID>95</GID>
<name>IN_1</name></connection>
<intersection>275.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>268.5,-33.5,268.5,-33</points>
<intersection>-33.5 2</intersection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>267.5,-33,268.5,-33</points>
<connection>
<GID>99</GID>
<name>OUT_0</name></connection>
<intersection>268.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>268.5,-33.5,269.5,-33.5</points>
<connection>
<GID>93</GID>
<name>IN_0</name></connection>
<intersection>268.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>268.5,-36,268.5,-35.5</points>
<intersection>-36 1</intersection>
<intersection>-35.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>267.5,-36,268.5,-36</points>
<connection>
<GID>101</GID>
<name>OUT_0</name></connection>
<intersection>268.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>268.5,-35.5,269.5,-35.5</points>
<connection>
<GID>93</GID>
<name>IN_1</name></connection>
<intersection>268.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>503.5,-38.5,523,-38.5</points>
<connection>
<GID>208</GID>
<name>IN_0</name></connection>
<connection>
<GID>216</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>282.5,-34.5,283.5,-34.5</points>
<connection>
<GID>95</GID>
<name>OUT</name></connection>
<connection>
<GID>115</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274.5,-45,274.5,-42.5</points>
<intersection>-45 2</intersection>
<intersection>-42.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>273.5,-42.5,274.5,-42.5</points>
<connection>
<GID>118</GID>
<name>OUT</name></connection>
<intersection>274.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>274.5,-45,275.5,-45</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>274.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274.5,-49.5,274.5,-47</points>
<intersection>-49.5 1</intersection>
<intersection>-47 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>273.5,-49.5,274.5,-49.5</points>
<connection>
<GID>119</GID>
<name>OUT</name></connection>
<intersection>274.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>274.5,-47,275.5,-47</points>
<connection>
<GID>120</GID>
<name>IN_1</name></connection>
<intersection>274.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>266.5,-43.5,266.5,-41.5</points>
<intersection>-43.5 3</intersection>
<intersection>-42.5 1</intersection>
<intersection>-41.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>266,-42.5,266.5,-42.5</points>
<connection>
<GID>121</GID>
<name>OUT_0</name></connection>
<intersection>266.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>266.5,-41.5,267.5,-41.5</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<intersection>266.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>266.5,-43.5,267.5,-43.5</points>
<connection>
<GID>118</GID>
<name>IN_1</name></connection>
<intersection>266.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>266.5,-50.5,266.5,-48.5</points>
<intersection>-50.5 3</intersection>
<intersection>-49.5 1</intersection>
<intersection>-48.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>266,-49.5,266.5,-49.5</points>
<connection>
<GID>122</GID>
<name>OUT_0</name></connection>
<intersection>266.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>266.5,-48.5,267.5,-48.5</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>266.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>266.5,-50.5,267.5,-50.5</points>
<connection>
<GID>119</GID>
<name>IN_1</name></connection>
<intersection>266.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>281.5,-46,282.5,-46</points>
<connection>
<GID>120</GID>
<name>OUT</name></connection>
<connection>
<GID>127</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274.5,-59.5,274.5,-57</points>
<intersection>-59.5 2</intersection>
<intersection>-57 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>273.5,-57,274.5,-57</points>
<connection>
<GID>144</GID>
<name>OUT</name></connection>
<intersection>274.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>274.5,-59.5,275.5,-59.5</points>
<connection>
<GID>149</GID>
<name>IN_0</name></connection>
<intersection>274.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>274.5,-64,274.5,-61.5</points>
<intersection>-64 1</intersection>
<intersection>-61.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>273.5,-64,274.5,-64</points>
<connection>
<GID>146</GID>
<name>OUT</name></connection>
<intersection>274.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>274.5,-61.5,275.5,-61.5</points>
<connection>
<GID>149</GID>
<name>IN_1</name></connection>
<intersection>274.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>266.5,-58,266.5,-56</points>
<intersection>-58 3</intersection>
<intersection>-57 1</intersection>
<intersection>-56 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>266,-57,266.5,-57</points>
<connection>
<GID>150</GID>
<name>OUT_0</name></connection>
<intersection>266.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>266.5,-56,267.5,-56</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<intersection>266.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>266.5,-58,267.5,-58</points>
<connection>
<GID>144</GID>
<name>IN_1</name></connection>
<intersection>266.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>266.5,-65,266.5,-63</points>
<intersection>-65 3</intersection>
<intersection>-64 1</intersection>
<intersection>-63 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>266,-64,266.5,-64</points>
<connection>
<GID>153</GID>
<name>OUT_0</name></connection>
<intersection>266.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>266.5,-63,267.5,-63</points>
<connection>
<GID>146</GID>
<name>IN_0</name></connection>
<intersection>266.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>266.5,-65,267.5,-65</points>
<connection>
<GID>146</GID>
<name>IN_1</name></connection>
<intersection>266.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>289,-60.5,290,-60.5</points>
<connection>
<GID>157</GID>
<name>OUT</name></connection>
<connection>
<GID>158</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>282,-61.5,282,-59.5</points>
<intersection>-61.5 3</intersection>
<intersection>-60.5 1</intersection>
<intersection>-59.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>281.5,-60.5,282,-60.5</points>
<connection>
<GID>149</GID>
<name>OUT</name></connection>
<intersection>282 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>282,-59.5,283,-59.5</points>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<intersection>282 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>282,-61.5,283,-61.5</points>
<connection>
<GID>157</GID>
<name>IN_1</name></connection>
<intersection>282 0</intersection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>285.5,-76.5,285.5,-74</points>
<intersection>-76.5 2</intersection>
<intersection>-74 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>284.5,-74,285.5,-74</points>
<connection>
<GID>160</GID>
<name>OUT</name></connection>
<intersection>285.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>285.5,-76.5,286.5,-76.5</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<intersection>285.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>285.5,-81,285.5,-78.5</points>
<intersection>-81 1</intersection>
<intersection>-78.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>284.5,-81,285.5,-81</points>
<connection>
<GID>161</GID>
<name>OUT</name></connection>
<intersection>285.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>285.5,-78.5,286.5,-78.5</points>
<connection>
<GID>162</GID>
<name>IN_1</name></connection>
<intersection>285.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>499.5,-53.5,499.5,-32.5</points>
<connection>
<GID>216</GID>
<name>IN_0</name></connection>
<connection>
<GID>199</GID>
<name>OUT_0</name></connection>
<intersection>-53.5 4</intersection>
<intersection>-46.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>499.5,-46.5,523,-46.5</points>
<connection>
<GID>212</GID>
<name>IN_0</name></connection>
<intersection>499.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>499.5,-53.5,523,-53.5</points>
<connection>
<GID>230</GID>
<name>IN_0</name></connection>
<intersection>499.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>509.5,-55.5,509.5,-32.5</points>
<connection>
<GID>219</GID>
<name>IN_0</name></connection>
<connection>
<GID>203</GID>
<name>OUT_0</name></connection>
<intersection>-55.5 4</intersection>
<intersection>-40.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>509.5,-40.5,523,-40.5</points>
<connection>
<GID>208</GID>
<name>IN_1</name></connection>
<intersection>509.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>509.5,-55.5,523,-55.5</points>
<connection>
<GID>230</GID>
<name>IN_1</name></connection>
<intersection>509.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>293,-78.5,293,-76.5</points>
<intersection>-78.5 3</intersection>
<intersection>-77.5 1</intersection>
<intersection>-76.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>292.5,-77.5,293,-77.5</points>
<connection>
<GID>162</GID>
<name>OUT</name></connection>
<intersection>293 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>293,-76.5,294,-76.5</points>
<connection>
<GID>163</GID>
<name>IN_0</name></connection>
<intersection>293 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>293,-78.5,294,-78.5</points>
<connection>
<GID>163</GID>
<name>IN_1</name></connection>
<intersection>293 0</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<hsegment>
<ID>9</ID>
<points>513.5,-48.5,523,-48.5</points>
<connection>
<GID>212</GID>
<name>IN_1</name></connection>
<connection>
<GID>219</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>277,-80,277,-75</points>
<intersection>-80 3</intersection>
<intersection>-77.5 1</intersection>
<intersection>-75 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>275.5,-77.5,277,-77.5</points>
<connection>
<GID>164</GID>
<name>OUT</name></connection>
<intersection>277 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>277,-75,278.5,-75</points>
<connection>
<GID>160</GID>
<name>IN_1</name></connection>
<intersection>277 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>277,-80,278.5,-80</points>
<connection>
<GID>161</GID>
<name>IN_0</name></connection>
<intersection>277 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>530,-42.5,530,-39.5</points>
<intersection>-42.5 1</intersection>
<intersection>-39.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>530,-42.5,531.5,-42.5</points>
<connection>
<GID>221</GID>
<name>IN_0</name></connection>
<intersection>530 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>529,-39.5,530,-39.5</points>
<connection>
<GID>208</GID>
<name>OUT</name></connection>
<intersection>530 0</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>265.5,-73,278.5,-73</points>
<connection>
<GID>160</GID>
<name>IN_0</name></connection>
<connection>
<GID>166</GID>
<name>OUT_0</name></connection>
<intersection>270 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>270,-76.5,270,-73</points>
<intersection>-76.5 5</intersection>
<intersection>-73 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>269.5,-76.5,270,-76.5</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<intersection>270 3</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>265.5,-82,278.5,-82</points>
<connection>
<GID>161</GID>
<name>IN_1</name></connection>
<connection>
<GID>167</GID>
<name>OUT_0</name></connection>
<intersection>270 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>270,-82,270,-78.5</points>
<intersection>-82 1</intersection>
<intersection>-78.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>269.5,-78.5,270,-78.5</points>
<connection>
<GID>164</GID>
<name>IN_1</name></connection>
<intersection>270 3</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>300,-77.5,301.5,-77.5</points>
<connection>
<GID>163</GID>
<name>OUT</name></connection>
<connection>
<GID>169</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>285.5,-93,285.5,-90.5</points>
<intersection>-93 2</intersection>
<intersection>-90.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>284.5,-90.5,285.5,-90.5</points>
<connection>
<GID>173</GID>
<name>OUT</name></connection>
<intersection>285.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>285.5,-93,286.5,-93</points>
<connection>
<GID>175</GID>
<name>IN_0</name></connection>
<intersection>285.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>285.5,-97.5,285.5,-95</points>
<intersection>-97.5 1</intersection>
<intersection>-95 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>284.5,-97.5,285.5,-97.5</points>
<connection>
<GID>174</GID>
<name>OUT</name></connection>
<intersection>285.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>285.5,-95,286.5,-95</points>
<connection>
<GID>175</GID>
<name>IN_1</name></connection>
<intersection>285.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>277,-96.5,277,-91.5</points>
<intersection>-96.5 3</intersection>
<intersection>-94 1</intersection>
<intersection>-91.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>275.5,-94,277,-94</points>
<connection>
<GID>176</GID>
<name>OUT</name></connection>
<intersection>277 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>277,-91.5,278.5,-91.5</points>
<connection>
<GID>173</GID>
<name>IN_1</name></connection>
<intersection>277 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>277,-96.5,278.5,-96.5</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<intersection>277 0</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>265.5,-89.5,278.5,-89.5</points>
<connection>
<GID>173</GID>
<name>IN_0</name></connection>
<connection>
<GID>177</GID>
<name>OUT_0</name></connection>
<intersection>270 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>270,-93,270,-89.5</points>
<intersection>-93 8</intersection>
<intersection>-89.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>269.5,-93,270,-93</points>
<connection>
<GID>176</GID>
<name>IN_0</name></connection>
<intersection>270 3</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>265.5,-98.5,278.5,-98.5</points>
<connection>
<GID>174</GID>
<name>IN_1</name></connection>
<connection>
<GID>178</GID>
<name>OUT_0</name></connection>
<intersection>270 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>270,-98.5,270,-95</points>
<intersection>-98.5 1</intersection>
<intersection>-95 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>269.5,-95,270,-95</points>
<connection>
<GID>176</GID>
<name>IN_1</name></connection>
<intersection>270 3</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>292.5,-94,294,-94</points>
<connection>
<GID>175</GID>
<name>OUT</name></connection>
<connection>
<GID>182</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>432,-40,432,-37.5</points>
<intersection>-40 2</intersection>
<intersection>-37.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>429,-37.5,432,-37.5</points>
<connection>
<GID>196</GID>
<name>OUT</name></connection>
<intersection>432 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>432,-40,435,-40</points>
<connection>
<GID>200</GID>
<name>IN_0</name></connection>
<intersection>432 0</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>432,-43.5,432,-42</points>
<intersection>-43.5 1</intersection>
<intersection>-42 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>429,-43.5,432,-43.5</points>
<connection>
<GID>198</GID>
<name>OUT</name></connection>
<intersection>432 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>432,-42,435,-42</points>
<connection>
<GID>200</GID>
<name>IN_1</name></connection>
<intersection>432 0</intersection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>364.5,-49.5,364.5,-32.5</points>
<connection>
<GID>202</GID>
<name>IN_0</name></connection>
<connection>
<GID>192</GID>
<name>OUT_0</name></connection>
<intersection>-49.5 11</intersection>
<intersection>-42.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>364.5,-42.5,423,-42.5</points>
<connection>
<GID>198</GID>
<name>IN_0</name></connection>
<intersection>364.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>364.5,-49.5,423,-49.5</points>
<connection>
<GID>205</GID>
<name>IN_0</name></connection>
<intersection>364.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>368.5,-36.5,423,-36.5</points>
<connection>
<GID>196</GID>
<name>IN_0</name></connection>
<connection>
<GID>202</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>375,-51.5,375,-32.5</points>
<connection>
<GID>204</GID>
<name>IN_0</name></connection>
<connection>
<GID>194</GID>
<name>OUT_0</name></connection>
<intersection>-51.5 7</intersection>
<intersection>-38.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>375,-38.5,423,-38.5</points>
<connection>
<GID>196</GID>
<name>IN_1</name></connection>
<intersection>375 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>375,-51.5,423,-51.5</points>
<connection>
<GID>205</GID>
<name>IN_1</name></connection>
<intersection>375 0</intersection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>379,-44.5,423,-44.5</points>
<connection>
<GID>198</GID>
<name>IN_1</name></connection>
<connection>
<GID>204</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>429,-50.5,432,-50.5</points>
<connection>
<GID>205</GID>
<name>OUT</name></connection>
<connection>
<GID>207</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>441,-41,442.5,-41</points>
<connection>
<GID>200</GID>
<name>OUT</name></connection>
<connection>
<GID>209</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>530,-47.5,530,-44.5</points>
<intersection>-47.5 2</intersection>
<intersection>-44.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>530,-44.5,531.5,-44.5</points>
<connection>
<GID>221</GID>
<name>IN_1</name></connection>
<intersection>530 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>529,-47.5,530,-47.5</points>
<connection>
<GID>212</GID>
<name>OUT</name></connection>
<intersection>530 0</intersection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>537.5,-43.5,539.5,-43.5</points>
<connection>
<GID>221</GID>
<name>OUT</name></connection>
<connection>
<GID>223</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>530,-55.5,530,-53.5</points>
<intersection>-55.5 3</intersection>
<intersection>-54.5 2</intersection>
<intersection>-53.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>530,-53.5,531,-53.5</points>
<connection>
<GID>232</GID>
<name>IN_0</name></connection>
<intersection>530 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>529,-54.5,530,-54.5</points>
<connection>
<GID>230</GID>
<name>OUT</name></connection>
<intersection>530 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>530,-55.5,531,-55.5</points>
<connection>
<GID>232</GID>
<name>IN_1</name></connection>
<intersection>530 0</intersection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>537,-54.5,539,-54.5</points>
<connection>
<GID>231</GID>
<name>N_in0</name></connection>
<connection>
<GID>232</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>616.5,-37.5,616.5,-26.5</points>
<connection>
<GID>246</GID>
<name>IN_0</name></connection>
<connection>
<GID>236</GID>
<name>OUT_0</name></connection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>616.5,-30.5,647.5,-30.5</points>
<connection>
<GID>240</GID>
<name>IN_0</name></connection>
<intersection>616.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>628.5,-39.5,628.5,-26.5</points>
<connection>
<GID>244</GID>
<name>IN_0</name></connection>
<connection>
<GID>238</GID>
<name>OUT_0</name></connection>
<intersection>-39.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>628.5,-39.5,647.5,-39.5</points>
<connection>
<GID>242</GID>
<name>IN_1</name></connection>
<intersection>628.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>632.5,-32.5,647.5,-32.5</points>
<connection>
<GID>240</GID>
<name>IN_1</name></connection>
<connection>
<GID>244</GID>
<name>OUT_0</name></connection>
<intersection>632.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>632.5,-44,632.5,-32.5</points>
<intersection>-44 4</intersection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>632.5,-44,648,-44</points>
<connection>
<GID>254</GID>
<name>IN_0</name></connection>
<intersection>632.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>620.5,-37.5,647.5,-37.5</points>
<connection>
<GID>242</GID>
<name>IN_0</name></connection>
<connection>
<GID>246</GID>
<name>OUT_0</name></connection>
<intersection>620.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>620.5,-46,620.5,-37.5</points>
<intersection>-46 4</intersection>
<intersection>-37.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>620.5,-46,648,-46</points>
<connection>
<GID>254</GID>
<name>IN_1</name></connection>
<intersection>620.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>655.5,-34,655.5,-31.5</points>
<intersection>-34 2</intersection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>653.5,-31.5,655.5,-31.5</points>
<connection>
<GID>240</GID>
<name>OUT</name></connection>
<intersection>655.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>655.5,-34,657.5,-34</points>
<connection>
<GID>248</GID>
<name>IN_0</name></connection>
<intersection>655.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>655.5,-38.5,655.5,-36</points>
<intersection>-38.5 1</intersection>
<intersection>-36 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>653.5,-38.5,655.5,-38.5</points>
<connection>
<GID>242</GID>
<name>OUT</name></connection>
<intersection>655.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>655.5,-36,657.5,-36</points>
<connection>
<GID>248</GID>
<name>IN_1</name></connection>
<intersection>655.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>664.5,-36,664.5,-34</points>
<intersection>-36 3</intersection>
<intersection>-35 1</intersection>
<intersection>-34 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>663.5,-35,664.5,-35</points>
<connection>
<GID>248</GID>
<name>OUT</name></connection>
<intersection>664.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>664.5,-34,666,-34</points>
<connection>
<GID>250</GID>
<name>IN_0</name></connection>
<intersection>664.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>664.5,-36,666,-36</points>
<connection>
<GID>250</GID>
<name>IN_1</name></connection>
<intersection>664.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>672,-35,674,-35</points>
<connection>
<GID>252</GID>
<name>N_in0</name></connection>
<connection>
<GID>250</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>655,-46,655,-44</points>
<intersection>-46 3</intersection>
<intersection>-45 1</intersection>
<intersection>-44 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>654,-45,655,-45</points>
<connection>
<GID>254</GID>
<name>OUT</name></connection>
<intersection>655 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>655,-44,656.5,-44</points>
<connection>
<GID>256</GID>
<name>IN_0</name></connection>
<intersection>655 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>655,-46,656.5,-46</points>
<connection>
<GID>256</GID>
<name>IN_1</name></connection>
<intersection>655 0</intersection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>662.5,-45,665,-45</points>
<connection>
<GID>258</GID>
<name>N_in0</name></connection>
<connection>
<GID>256</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>-0.00025201,33.5808,338.954,-133.958</PageViewport></page 2>
<page 3>
<PageViewport>-0.00025201,33.5808,338.954,-133.958</PageViewport></page 3>
<page 4>
<PageViewport>-0.00025201,33.5808,338.954,-133.958</PageViewport></page 4>
<page 5>
<PageViewport>-0.00025201,33.5808,338.954,-133.958</PageViewport></page 5>
<page 6>
<PageViewport>-0.00025201,33.5808,338.954,-133.958</PageViewport></page 6>
<page 7>
<PageViewport>-0.00025201,33.5808,338.954,-133.958</PageViewport></page 7>
<page 8>
<PageViewport>-0.00025201,33.5808,338.954,-133.958</PageViewport></page 8>
<page 9>
<PageViewport>-0.00025201,33.5808,338.954,-133.958</PageViewport></page 9></circuit>