<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-9,6,113.4,-54.5</PageViewport>
<gate>
<ID>2</ID>
<type>AA_MUX_2x1</type>
<position>13,-17</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>3 </output>
<input>
<ID>SEL_0</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_LABEL</type>
<position>12.5,-5</position>
<gparam>LABEL_TEXT 2*1 MUX</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>4,-14</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>3.5,-18</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>10</ID>
<type>GA_LED</type>
<position>19,-17</position>
<input>
<ID>N_in0</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>10,-9.5</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>14</ID>
<type>AE_MUX_4x1</type>
<position>48.5,-14.5</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>7 </input>
<input>
<ID>IN_2</ID>6 </input>
<input>
<ID>IN_3</ID>5 </input>
<output>
<ID>OUT</ID>9 </output>
<input>
<ID>SEL_0</ID>23 </input>
<input>
<ID>SEL_1</ID>22 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_TOGGLE</type>
<position>39.5,-11</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_TOGGLE</type>
<position>39.5,-14</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_TOGGLE</type>
<position>39.5,-16.5</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_TOGGLE</type>
<position>39.5,-19</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>24</ID>
<type>GA_LED</type>
<position>56.5,-14.5</position>
<input>
<ID>N_in0</ID>9 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>AI_MUX_8x1</type>
<position>84.5,-14.5</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>16 </input>
<input>
<ID>IN_2</ID>15 </input>
<input>
<ID>IN_3</ID>14 </input>
<input>
<ID>IN_4</ID>13 </input>
<input>
<ID>IN_5</ID>12 </input>
<input>
<ID>IN_6</ID>11 </input>
<input>
<ID>IN_7</ID>10 </input>
<output>
<ID>OUT</ID>21 </output>
<input>
<ID>SEL_0</ID>19 </input>
<input>
<ID>SEL_1</ID>20 </input>
<input>
<ID>SEL_2</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_TOGGLE</type>
<position>72,-9</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_TOGGLE</type>
<position>72,-12.5</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>34</ID>
<type>AA_TOGGLE</type>
<position>72,-15.5</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_TOGGLE</type>
<position>72,-19.5</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_TOGGLE</type>
<position>72,-23.5</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>40</ID>
<type>AA_TOGGLE</type>
<position>72,-27.5</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_TOGGLE</type>
<position>80,-6.5</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_TOGGLE</type>
<position>81,-29.5</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_TOGGLE</type>
<position>44.5,-5.5</position>
<output>
<ID>OUT_0</ID>22 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>48</ID>
<type>AA_TOGGLE</type>
<position>50.5,-5</position>
<output>
<ID>OUT_0</ID>23 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_TOGGLE</type>
<position>83,-4.5</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>52</ID>
<type>AA_TOGGLE</type>
<position>85.5,-4.5</position>
<output>
<ID>OUT_0</ID>20 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>54</ID>
<type>AA_TOGGLE</type>
<position>88,-4.5</position>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>56</ID>
<type>GA_LED</type>
<position>93,-14</position>
<input>
<ID>N_in0</ID>21 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>58</ID>
<type>AA_LABEL</type>
<position>-3,-13.5</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>60</ID>
<type>AA_LABEL</type>
<position>-2.5,-17.5</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>61</ID>
<type>AA_LABEL</type>
<position>34.5,-11</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>62</ID>
<type>AA_LABEL</type>
<position>77,-5.5</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>63</ID>
<type>AA_LABEL</type>
<position>35,-13.5</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>64</ID>
<type>AA_LABEL</type>
<position>68,-9.5</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>66</ID>
<type>AA_LABEL</type>
<position>35,-16.5</position>
<gparam>LABEL_TEXT D2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>AA_LABEL</type>
<position>35,-19</position>
<gparam>LABEL_TEXT D3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>69</ID>
<type>AA_LABEL</type>
<position>68.5,-15</position>
<gparam>LABEL_TEXT D3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>AA_LABEL</type>
<position>68,-12</position>
<gparam>LABEL_TEXT D2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>72</ID>
<type>AA_LABEL</type>
<position>68.5,-19</position>
<gparam>LABEL_TEXT D4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>74</ID>
<type>AA_LABEL</type>
<position>68.5,-23.5</position>
<gparam>LABEL_TEXT D5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>76</ID>
<type>AA_LABEL</type>
<position>68.5,-27.5</position>
<gparam>LABEL_TEXT D6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>78</ID>
<type>AA_LABEL</type>
<position>81,-32.5</position>
<gparam>LABEL_TEXT D7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>80</ID>
<type>AA_LABEL</type>
<position>13,-9</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>82</ID>
<type>AA_LABEL</type>
<position>50.5,-2.5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>84</ID>
<type>AA_LABEL</type>
<position>88.5,-2</position>
<gparam>LABEL_TEXT S2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>86</ID>
<type>AA_LABEL</type>
<position>86,2</position>
<gparam>LABEL_TEXT 8*1 MUX</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>87</ID>
<type>AA_LABEL</type>
<position>44,-3</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>88</ID>
<type>AA_LABEL</type>
<position>82,-2</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>89</ID>
<type>AA_LABEL</type>
<position>85.5,-2</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>91</ID>
<type>AA_LABEL</type>
<position>47,1.5</position>
<gparam>LABEL_TEXT 4*1 MUX</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-16,9,-14</points>
<intersection>-16 1</intersection>
<intersection>-14 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-16,11,-16</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>9 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>6,-14,9,-14</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>9 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5.5,-18,11,-18</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>15,-17,18,-17</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<connection>
<GID>10</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10,-14.5,10,-11.5</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>10,-14.5,13,-14.5</points>
<connection>
<GID>2</GID>
<name>SEL_0</name></connection>
<intersection>10 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-11.5,43.5,-11</points>
<intersection>-11.5 1</intersection>
<intersection>-11 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43.5,-11.5,45.5,-11.5</points>
<connection>
<GID>14</GID>
<name>IN_3</name></connection>
<intersection>43.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>41.5,-11,43.5,-11</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-14,43.5,-13.5</points>
<intersection>-14 2</intersection>
<intersection>-13.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43.5,-13.5,45.5,-13.5</points>
<connection>
<GID>14</GID>
<name>IN_2</name></connection>
<intersection>43.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>41.5,-14,43.5,-14</points>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-16.5,43.5,-15.5</points>
<intersection>-16.5 2</intersection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43.5,-15.5,45.5,-15.5</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>43.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>41.5,-16.5,43.5,-16.5</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-19,43.5,-17.5</points>
<intersection>-19 2</intersection>
<intersection>-17.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43.5,-17.5,45.5,-17.5</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>43.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>41.5,-19,43.5,-19</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>51.5,-14.5,55.5,-14.5</points>
<connection>
<GID>24</GID>
<name>N_in0</name></connection>
<connection>
<GID>14</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-11,80,-8.5</points>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80,-11,81.5,-11</points>
<connection>
<GID>28</GID>
<name>IN_7</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79.5,-12,79.5,-9</points>
<intersection>-12 1</intersection>
<intersection>-9 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>79.5,-12,81.5,-12</points>
<connection>
<GID>28</GID>
<name>IN_6</name></connection>
<intersection>79.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>74,-9,79.5,-9</points>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection>
<intersection>79.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79.5,-13,79.5,-12.5</points>
<intersection>-13 1</intersection>
<intersection>-12.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>79.5,-13,81.5,-13</points>
<connection>
<GID>28</GID>
<name>IN_5</name></connection>
<intersection>79.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>74,-12.5,79.5,-12.5</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<intersection>79.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74,-14.5,81.5,-14.5</points>
<intersection>74 5</intersection>
<intersection>81.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>81.5,-14.5,81.5,-14</points>
<connection>
<GID>28</GID>
<name>IN_4</name></connection>
<intersection>-14.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>74,-15.5,74,-14.5</points>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78,-19.5,78,-15</points>
<intersection>-19.5 2</intersection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>78,-15,81.5,-15</points>
<connection>
<GID>28</GID>
<name>IN_3</name></connection>
<intersection>78 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>74,-19.5,78,-19.5</points>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<intersection>78 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79,-23.5,79,-16</points>
<intersection>-23.5 2</intersection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>79,-16,81.5,-16</points>
<connection>
<GID>28</GID>
<name>IN_2</name></connection>
<intersection>79 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>74,-23.5,79,-23.5</points>
<connection>
<GID>38</GID>
<name>OUT_0</name></connection>
<intersection>79 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79.5,-27.5,79.5,-17</points>
<intersection>-27.5 2</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>79.5,-17,81.5,-17</points>
<connection>
<GID>28</GID>
<name>IN_1</name></connection>
<intersection>79.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>74,-27.5,79.5,-27.5</points>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection>
<intersection>79.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,-27.5,81,-18</points>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>81,-18,81.5,-18</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>81 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83,-7.5,83,-6.5</points>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection>
<intersection>-7.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>83.5,-9,83.5,-7.5</points>
<connection>
<GID>28</GID>
<name>SEL_2</name></connection>
<intersection>-7.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>83,-7.5,83.5,-7.5</points>
<intersection>83 0</intersection>
<intersection>83.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,-7.5,88,-6.5</points>
<connection>
<GID>54</GID>
<name>OUT_0</name></connection>
<intersection>-7.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>85.5,-9,85.5,-7.5</points>
<connection>
<GID>28</GID>
<name>SEL_0</name></connection>
<intersection>-7.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>85.5,-7.5,88,-7.5</points>
<intersection>85.5 1</intersection>
<intersection>88 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85.5,-7,85.5,-6.5</points>
<connection>
<GID>52</GID>
<name>OUT_0</name></connection>
<intersection>-7 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>84.5,-9,84.5,-7</points>
<connection>
<GID>28</GID>
<name>SEL_1</name></connection>
<intersection>-7 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>84.5,-7,85.5,-7</points>
<intersection>84.5 1</intersection>
<intersection>85.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-14.5,89.5,-14</points>
<intersection>-14.5 2</intersection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>89.5,-14,92,-14</points>
<connection>
<GID>56</GID>
<name>N_in0</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>87.5,-14.5,89.5,-14.5</points>
<connection>
<GID>28</GID>
<name>OUT</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48.5,-9.5,48.5,-5.5</points>
<connection>
<GID>14</GID>
<name>SEL_1</name></connection>
<intersection>-5.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46.5,-5.5,48.5,-5.5</points>
<connection>
<GID>46</GID>
<name>OUT_0</name></connection>
<intersection>48.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-9.5,49.5,-8</points>
<connection>
<GID>14</GID>
<name>SEL_0</name></connection>
<intersection>-8 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>50.5,-8,50.5,-7</points>
<connection>
<GID>48</GID>
<name>OUT_0</name></connection>
<intersection>-8 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>49.5,-8,50.5,-8</points>
<intersection>49.5 0</intersection>
<intersection>50.5 1</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-19.5257,5.26646,69.5257,-38.75</PageViewport>
<gate>
<ID>93</ID>
<type>AA_MUX_2x1</type>
<position>17.5,-10</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>30 </input>
<output>
<ID>OUT</ID>26 </output>
<input>
<ID>SEL_0</ID>41 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>95</ID>
<type>AA_MUX_2x1</type>
<position>17.5,-18</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>27 </output>
<input>
<ID>SEL_0</ID>41 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>97</ID>
<type>AA_MUX_2x1</type>
<position>17.5,-26.5</position>
<input>
<ID>IN_0</ID>35 </input>
<input>
<ID>IN_1</ID>34 </input>
<output>
<ID>OUT</ID>28 </output>
<input>
<ID>SEL_0</ID>41 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>99</ID>
<type>AA_MUX_2x1</type>
<position>17.5,-34.5</position>
<input>
<ID>IN_0</ID>37 </input>
<input>
<ID>IN_1</ID>36 </input>
<output>
<ID>OUT</ID>29 </output>
<input>
<ID>SEL_0</ID>41 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>101</ID>
<type>AA_MUX_2x1</type>
<position>27.5,-13.5</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>24 </output>
<input>
<ID>SEL_0</ID>40 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>103</ID>
<type>AA_MUX_2x1</type>
<position>28,-29.5</position>
<input>
<ID>IN_0</ID>29 </input>
<input>
<ID>IN_1</ID>28 </input>
<output>
<ID>OUT</ID>25 </output>
<input>
<ID>SEL_0</ID>40 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>105</ID>
<type>AA_MUX_2x1</type>
<position>37.5,-21</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>38 </output>
<input>
<ID>SEL_0</ID>43 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>107</ID>
<type>AA_TOGGLE</type>
<position>5.5,-9</position>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>109</ID>
<type>AA_TOGGLE</type>
<position>5,-13</position>
<output>
<ID>OUT_0</ID>31 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>111</ID>
<type>AA_TOGGLE</type>
<position>5,-16.5</position>
<output>
<ID>OUT_0</ID>32 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>113</ID>
<type>AA_TOGGLE</type>
<position>4.5,-20</position>
<output>
<ID>OUT_0</ID>33 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>115</ID>
<type>AA_TOGGLE</type>
<position>5,-25</position>
<output>
<ID>OUT_0</ID>34 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>117</ID>
<type>AA_TOGGLE</type>
<position>4.5,-29</position>
<output>
<ID>OUT_0</ID>35 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>119</ID>
<type>AA_TOGGLE</type>
<position>5,-33</position>
<output>
<ID>OUT_0</ID>36 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>121</ID>
<type>AA_TOGGLE</type>
<position>5,-37.5</position>
<output>
<ID>OUT_0</ID>37 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>123</ID>
<type>GA_LED</type>
<position>49,-21</position>
<input>
<ID>N_in0</ID>38 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>125</ID>
<type>AA_LABEL</type>
<position>1.5,-37.5</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>126</ID>
<type>AA_LABEL</type>
<position>1.5,-33</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>127</ID>
<type>AA_LABEL</type>
<position>1,-29</position>
<gparam>LABEL_TEXT D2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>128</ID>
<type>AA_LABEL</type>
<position>1.5,-24.5</position>
<gparam>LABEL_TEXT D3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>129</ID>
<type>AA_LABEL</type>
<position>1.5,-19.5</position>
<gparam>LABEL_TEXT D4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>130</ID>
<type>AA_LABEL</type>
<position>1,-16</position>
<gparam>LABEL_TEXT D5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>131</ID>
<type>AA_LABEL</type>
<position>1.5,-12.5</position>
<gparam>LABEL_TEXT D6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>132</ID>
<type>AA_LABEL</type>
<position>2,-9</position>
<gparam>LABEL_TEXT D7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>134</ID>
<type>AA_TOGGLE</type>
<position>18,-1</position>
<output>
<ID>OUT_0</ID>41 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>136</ID>
<type>AA_TOGGLE</type>
<position>27.5,-5</position>
<output>
<ID>OUT_0</ID>40 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>138</ID>
<type>AA_TOGGLE</type>
<position>37,-11.5</position>
<output>
<ID>OUT_0</ID>43 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>139</ID>
<type>AA_LABEL</type>
<position>16.5,1</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>140</ID>
<type>AA_LABEL</type>
<position>27,-2</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>141</ID>
<type>AA_LABEL</type>
<position>37,-8.5</position>
<gparam>LABEL_TEXT S2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>143</ID>
<type>AA_LABEL</type>
<position>21.5,4.5</position>
<gparam>LABEL_TEXT 8*1 USING 2*1 MUX</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-20,32,-13.5</points>
<intersection>-20 1</intersection>
<intersection>-13.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,-20,35.5,-20</points>
<connection>
<GID>105</GID>
<name>IN_1</name></connection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29.5,-13.5,32,-13.5</points>
<connection>
<GID>101</GID>
<name>OUT</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-29.5,32.5,-22</points>
<intersection>-29.5 2</intersection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-22,35.5,-22</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30,-29.5,32.5,-29.5</points>
<connection>
<GID>103</GID>
<name>OUT</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-12.5,22.5,-10</points>
<intersection>-12.5 1</intersection>
<intersection>-10 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-12.5,25.5,-12.5</points>
<connection>
<GID>101</GID>
<name>IN_1</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>19.5,-10,22.5,-10</points>
<connection>
<GID>93</GID>
<name>OUT</name></connection>
<intersection>22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-18,22,-14.5</points>
<intersection>-18 2</intersection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22,-14.5,25.5,-14.5</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>22 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>19.5,-18,22,-18</points>
<connection>
<GID>95</GID>
<name>OUT</name></connection>
<intersection>22 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-28.5,22.5,-26.5</points>
<intersection>-28.5 1</intersection>
<intersection>-26.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-28.5,26,-28.5</points>
<connection>
<GID>103</GID>
<name>IN_1</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>19.5,-26.5,22.5,-26.5</points>
<connection>
<GID>97</GID>
<name>OUT</name></connection>
<intersection>22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-34.5,22.5,-30.5</points>
<intersection>-34.5 2</intersection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-30.5,26,-30.5</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>19.5,-34.5,22.5,-34.5</points>
<connection>
<GID>99</GID>
<name>OUT</name></connection>
<intersection>22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7.5,-9,15.5,-9</points>
<connection>
<GID>93</GID>
<name>IN_1</name></connection>
<connection>
<GID>107</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>9,-11,15.5,-11</points>
<connection>
<GID>93</GID>
<name>IN_0</name></connection>
<intersection>9 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>9,-13,9,-11</points>
<intersection>-13 4</intersection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>7,-13,9,-13</points>
<connection>
<GID>109</GID>
<name>OUT_0</name></connection>
<intersection>9 3</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12.5,-17,12.5,-16.5</points>
<intersection>-17 1</intersection>
<intersection>-16.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>12.5,-17,15.5,-17</points>
<connection>
<GID>95</GID>
<name>IN_1</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>7,-16.5,12.5,-16.5</points>
<connection>
<GID>111</GID>
<name>OUT_0</name></connection>
<intersection>12.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12.5,-20,12.5,-19</points>
<intersection>-20 2</intersection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>12.5,-19,15.5,-19</points>
<connection>
<GID>95</GID>
<name>IN_0</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>6.5,-20,12.5,-20</points>
<connection>
<GID>113</GID>
<name>OUT_0</name></connection>
<intersection>12.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12.5,-25.5,12.5,-25</points>
<intersection>-25.5 1</intersection>
<intersection>-25 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>12.5,-25.5,15.5,-25.5</points>
<connection>
<GID>97</GID>
<name>IN_1</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>7,-25,12.5,-25</points>
<connection>
<GID>115</GID>
<name>OUT_0</name></connection>
<intersection>12.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6.5,-29,15.5,-29</points>
<connection>
<GID>117</GID>
<name>OUT_0</name></connection>
<intersection>15.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>15.5,-29,15.5,-27.5</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<intersection>-29 1</intersection></vsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12.5,-33.5,12.5,-33</points>
<intersection>-33.5 1</intersection>
<intersection>-33 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>12.5,-33.5,15.5,-33.5</points>
<connection>
<GID>99</GID>
<name>IN_1</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>7,-33,12.5,-33</points>
<connection>
<GID>119</GID>
<name>OUT_0</name></connection>
<intersection>12.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12.5,-37.5,12.5,-35.5</points>
<intersection>-37.5 2</intersection>
<intersection>-35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>12.5,-35.5,15.5,-35.5</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>7,-37.5,12.5,-37.5</points>
<connection>
<GID>121</GID>
<name>OUT_0</name></connection>
<intersection>12.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39.5,-21,48,-21</points>
<connection>
<GID>105</GID>
<name>OUT</name></connection>
<connection>
<GID>123</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-16.5,27.5,-7</points>
<connection>
<GID>136</GID>
<name>OUT_0</name></connection>
<connection>
<GID>101</GID>
<name>SEL_0</name></connection>
<intersection>-16.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>28,-27,28,-16.5</points>
<connection>
<GID>103</GID>
<name>SEL_0</name></connection>
<intersection>-16.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>27.5,-16.5,28,-16.5</points>
<intersection>27.5 0</intersection>
<intersection>28 1</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-32,17.5,-3</points>
<connection>
<GID>97</GID>
<name>SEL_0</name></connection>
<connection>
<GID>93</GID>
<name>SEL_0</name></connection>
<connection>
<GID>99</GID>
<name>SEL_0</name></connection>
<connection>
<GID>95</GID>
<name>SEL_0</name></connection>
<intersection>-3 24</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>17.5,-3,18,-3</points>
<connection>
<GID>134</GID>
<name>OUT_0</name></connection>
<intersection>17.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,-18.5,37.5,-13.5</points>
<connection>
<GID>105</GID>
<name>SEL_0</name></connection>
<intersection>-13.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>37,-13.5,37.5,-13.5</points>
<connection>
<GID>138</GID>
<name>OUT_0</name></connection>
<intersection>37.5 0</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>-36,0,86.4,-60.5</PageViewport>
<gate>
<ID>145</ID>
<type>AA_AND3</type>
<position>27,-13</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>49 </input>
<input>
<ID>IN_2</ID>44 </input>
<output>
<ID>OUT</ID>51 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>149</ID>
<type>AA_AND3</type>
<position>27.5,-30</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>46 </input>
<input>
<ID>IN_2</ID>44 </input>
<output>
<ID>OUT</ID>53 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>151</ID>
<type>AA_AND3</type>
<position>27.5,-38.5</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>IN_1</ID>46 </input>
<input>
<ID>IN_2</ID>44 </input>
<output>
<ID>OUT</ID>54 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>153</ID>
<type>AA_TOGGLE</type>
<position>-19.5,-17</position>
<output>
<ID>OUT_0</ID>45 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>155</ID>
<type>AA_TOGGLE</type>
<position>-20,-24</position>
<output>
<ID>OUT_0</ID>46 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>157</ID>
<type>AA_TOGGLE</type>
<position>-19.5,-40</position>
<output>
<ID>OUT_0</ID>44 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>161</ID>
<type>AE_SMALL_INVERTER</type>
<position>-5,-26.5</position>
<input>
<ID>IN_0</ID>46 </input>
<output>
<ID>OUT_0</ID>49 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>163</ID>
<type>AE_SMALL_INVERTER</type>
<position>-7.5,-13.5</position>
<input>
<ID>IN_0</ID>45 </input>
<output>
<ID>OUT_0</ID>50 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>165</ID>
<type>AA_LABEL</type>
<position>-28,-16</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>167</ID>
<type>AA_LABEL</type>
<position>-28,-23.5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>169</ID>
<type>AA_LABEL</type>
<position>-25,-39.5</position>
<gparam>LABEL_TEXT Din</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>171</ID>
<type>AA_LABEL</type>
<position>45,-12.5</position>
<gparam>LABEL_TEXT I0= Din S1' S0'</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>178</ID>
<type>AA_LABEL</type>
<position>44.5,-21</position>
<gparam>LABEL_TEXT I1= Din S1' S0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>179</ID>
<type>AA_LABEL</type>
<position>43.5,-29.5</position>
<gparam>LABEL_TEXT I2= Din S1 S0'</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>180</ID>
<type>AA_LABEL</type>
<position>43.5,-38.5</position>
<gparam>LABEL_TEXT I3= Din S1 S0</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>182</ID>
<type>AA_AND3</type>
<position>27.5,-21.5</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>IN_1</ID>49 </input>
<input>
<ID>IN_2</ID>44 </input>
<output>
<ID>OUT</ID>52 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>184</ID>
<type>GA_LED</type>
<position>31,-13</position>
<input>
<ID>N_in0</ID>51 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>186</ID>
<type>GA_LED</type>
<position>31.5,-21.5</position>
<input>
<ID>N_in0</ID>52 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>188</ID>
<type>GA_LED</type>
<position>31.5,-30</position>
<input>
<ID>N_in0</ID>53 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>190</ID>
<type>GA_LED</type>
<position>31.5,-38.5</position>
<input>
<ID>N_in0</ID>54 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>44</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-18,-40.5,24.5,-40.5</points>
<connection>
<GID>151</GID>
<name>IN_2</name></connection>
<intersection>-18 10</intersection>
<intersection>10.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>10.5,-40.5,10.5,-15</points>
<intersection>-40.5 1</intersection>
<intersection>-32 7</intersection>
<intersection>-23.5 12</intersection>
<intersection>-15 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>10.5,-15,24,-15</points>
<connection>
<GID>145</GID>
<name>IN_2</name></connection>
<intersection>10.5 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>10.5,-32,24.5,-32</points>
<connection>
<GID>149</GID>
<name>IN_2</name></connection>
<intersection>10.5 3</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-18,-40.5,-18,-40</points>
<intersection>-40.5 1</intersection>
<intersection>-40 13</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>10.5,-23.5,24.5,-23.5</points>
<connection>
<GID>182</GID>
<name>IN_2</name></connection>
<intersection>10.5 3</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-18,-40,-17.5,-40</points>
<connection>
<GID>157</GID>
<name>OUT_0</name></connection>
<intersection>-18 10</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-17.5,-17,-9.5,-17</points>
<connection>
<GID>153</GID>
<name>OUT_0</name></connection>
<intersection>-9.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-9.5,-36.5,-9.5,-13.5</points>
<connection>
<GID>163</GID>
<name>IN_0</name></connection>
<intersection>-36.5 7</intersection>
<intersection>-19.5 9</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-9.5,-36.5,24.5,-36.5</points>
<connection>
<GID>151</GID>
<name>IN_0</name></connection>
<intersection>-9.5 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-9.5,-19.5,24.5,-19.5</points>
<connection>
<GID>182</GID>
<name>IN_0</name></connection>
<intersection>-9.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-18,-21.5,-1.5,-21.5</points>
<intersection>-18 8</intersection>
<intersection>-7.5 5</intersection>
<intersection>-1.5 9</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-7.5,-26.5,-7.5,-21.5</points>
<intersection>-26.5 7</intersection>
<intersection>-21.5 2</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-7.5,-26.5,-7,-26.5</points>
<connection>
<GID>161</GID>
<name>IN_0</name></connection>
<intersection>-7.5 5</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-18,-24,-18,-21.5</points>
<connection>
<GID>155</GID>
<name>OUT_0</name></connection>
<intersection>-21.5 2</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>-1.5,-38.5,-1.5,-21.5</points>
<intersection>-38.5 12</intersection>
<intersection>-30 10</intersection>
<intersection>-21.5 2</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>-1.5,-30,24.5,-30</points>
<connection>
<GID>149</GID>
<name>IN_1</name></connection>
<intersection>-1.5 9</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-1.5,-38.5,24.5,-38.5</points>
<connection>
<GID>151</GID>
<name>IN_1</name></connection>
<intersection>-1.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9.5,-24.5,9.5,-13</points>
<intersection>-24.5 1</intersection>
<intersection>-21.5 5</intersection>
<intersection>-13 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-3,-24.5,9.5,-24.5</points>
<intersection>-3 3</intersection>
<intersection>9.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>9.5,-13,24,-13</points>
<connection>
<GID>145</GID>
<name>IN_1</name></connection>
<intersection>9.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-3,-26.5,-3,-24.5</points>
<connection>
<GID>161</GID>
<name>OUT_0</name></connection>
<intersection>-24.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>9.5,-21.5,24.5,-21.5</points>
<connection>
<GID>182</GID>
<name>IN_1</name></connection>
<intersection>9.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4,-28,4,-11</points>
<intersection>-28 4</intersection>
<intersection>-13.5 2</intersection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>4,-11,24,-11</points>
<connection>
<GID>145</GID>
<name>IN_0</name></connection>
<intersection>4 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-5.5,-13.5,4,-13.5</points>
<connection>
<GID>163</GID>
<name>OUT_0</name></connection>
<intersection>4 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>4,-28,24.5,-28</points>
<connection>
<GID>149</GID>
<name>IN_0</name></connection>
<intersection>4 0</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-13,30,-13</points>
<connection>
<GID>184</GID>
<name>N_in0</name></connection>
<connection>
<GID>145</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-21.5,30.5,-21.5</points>
<connection>
<GID>186</GID>
<name>N_in0</name></connection>
<connection>
<GID>182</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-30,30.5,-30</points>
<connection>
<GID>188</GID>
<name>N_in0</name></connection>
<connection>
<GID>149</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-38.5,30.5,-38.5</points>
<connection>
<GID>190</GID>
<name>N_in0</name></connection>
<connection>
<GID>151</GID>
<name>OUT</name></connection></vsegment></shape></wire></page 2>
<page 3>
<PageViewport>-47.0667,12.8667,116.133,-67.8</PageViewport>
<gate>
<ID>194</ID>
<type>AA_AND4</type>
<position>44,-8.5</position>
<input>
<ID>IN_0</ID>55 </input>
<input>
<ID>IN_1</ID>61 </input>
<input>
<ID>IN_2</ID>60 </input>
<input>
<ID>IN_3</ID>56 </input>
<output>
<ID>OUT</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>196</ID>
<type>AA_AND4</type>
<position>44,-17.5</position>
<input>
<ID>IN_0</ID>55 </input>
<input>
<ID>IN_1</ID>61 </input>
<input>
<ID>IN_2</ID>57 </input>
<input>
<ID>IN_3</ID>59 </input>
<output>
<ID>OUT</ID>64 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>198</ID>
<type>AA_AND4</type>
<position>44,-26.5</position>
<input>
<ID>IN_0</ID>55 </input>
<input>
<ID>IN_1</ID>61 </input>
<input>
<ID>IN_2</ID>57 </input>
<input>
<ID>IN_3</ID>56 </input>
<output>
<ID>OUT</ID>65 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>200</ID>
<type>AA_AND4</type>
<position>44,-35.5</position>
<input>
<ID>IN_0</ID>55 </input>
<input>
<ID>IN_1</ID>58 </input>
<input>
<ID>IN_2</ID>60 </input>
<input>
<ID>IN_3</ID>59 </input>
<output>
<ID>OUT</ID>66 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>202</ID>
<type>AA_AND4</type>
<position>44,-44.5</position>
<input>
<ID>IN_0</ID>55 </input>
<input>
<ID>IN_1</ID>58 </input>
<input>
<ID>IN_2</ID>60 </input>
<input>
<ID>IN_3</ID>56 </input>
<output>
<ID>OUT</ID>67 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>204</ID>
<type>AA_AND4</type>
<position>44,-53.5</position>
<input>
<ID>IN_0</ID>55 </input>
<input>
<ID>IN_1</ID>59 </input>
<input>
<ID>IN_2</ID>58 </input>
<input>
<ID>IN_3</ID>57 </input>
<output>
<ID>OUT</ID>68 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>206</ID>
<type>AA_AND4</type>
<position>44,-62.5</position>
<input>
<ID>IN_0</ID>55 </input>
<input>
<ID>IN_1</ID>58 </input>
<input>
<ID>IN_2</ID>57 </input>
<input>
<ID>IN_3</ID>56 </input>
<output>
<ID>OUT</ID>69 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>208</ID>
<type>AA_TOGGLE</type>
<position>-2,7.5</position>
<output>
<ID>OUT_0</ID>57 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>210</ID>
<type>AA_TOGGLE</type>
<position>6.5,7.5</position>
<output>
<ID>OUT_0</ID>58 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>212</ID>
<type>AA_TOGGLE</type>
<position>15.5,7.5</position>
<output>
<ID>OUT_0</ID>55 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>214</ID>
<type>AA_TOGGLE</type>
<position>-10.5,7.5</position>
<output>
<ID>OUT_0</ID>56 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>216</ID>
<type>AE_SMALL_INVERTER</type>
<position>-7,5</position>
<input>
<ID>IN_0</ID>56 </input>
<output>
<ID>OUT_0</ID>59 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>218</ID>
<type>AE_SMALL_INVERTER</type>
<position>2,5</position>
<input>
<ID>IN_0</ID>57 </input>
<output>
<ID>OUT_0</ID>60 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>220</ID>
<type>AE_SMALL_INVERTER</type>
<position>11,5</position>
<input>
<ID>IN_0</ID>58 </input>
<output>
<ID>OUT_0</ID>61 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>224</ID>
<type>GA_LED</type>
<position>48,0.5</position>
<input>
<ID>N_in0</ID>62 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>226</ID>
<type>GA_LED</type>
<position>48,-8.5</position>
<input>
<ID>N_in0</ID>63 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>228</ID>
<type>GA_LED</type>
<position>48,-17.5</position>
<input>
<ID>N_in0</ID>64 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>230</ID>
<type>GA_LED</type>
<position>48,-26.5</position>
<input>
<ID>N_in0</ID>65 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>232</ID>
<type>GA_LED</type>
<position>48,-35.5</position>
<input>
<ID>N_in0</ID>66 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>234</ID>
<type>GA_LED</type>
<position>48,-44.5</position>
<input>
<ID>N_in0</ID>67 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>236</ID>
<type>GA_LED</type>
<position>48,-53.5</position>
<input>
<ID>N_in0</ID>68 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>238</ID>
<type>GA_LED</type>
<position>48,-62.5</position>
<input>
<ID>N_in0</ID>69 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>240</ID>
<type>AA_LABEL</type>
<position>55,1</position>
<gparam>LABEL_TEXT I0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>241</ID>
<type>AA_LABEL</type>
<position>55.5,-8</position>
<gparam>LABEL_TEXT I1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>242</ID>
<type>AA_LABEL</type>
<position>55.5,-16.5</position>
<gparam>LABEL_TEXT I2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>243</ID>
<type>AA_LABEL</type>
<position>55,-26.5</position>
<gparam>LABEL_TEXT I3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>244</ID>
<type>AA_LABEL</type>
<position>55,-35.5</position>
<gparam>LABEL_TEXT I4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>245</ID>
<type>AA_LABEL</type>
<position>55,-44</position>
<gparam>LABEL_TEXT I5</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>246</ID>
<type>AA_LABEL</type>
<position>54.5,-53.5</position>
<gparam>LABEL_TEXT I6</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>247</ID>
<type>AA_LABEL</type>
<position>55,-61.5</position>
<gparam>LABEL_TEXT I7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>192</ID>
<type>AA_AND4</type>
<position>44,0.5</position>
<input>
<ID>IN_0</ID>55 </input>
<input>
<ID>IN_1</ID>61 </input>
<input>
<ID>IN_2</ID>60 </input>
<input>
<ID>IN_3</ID>59 </input>
<output>
<ID>OUT</ID>62 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15.5,-59.5,15.5,5.5</points>
<connection>
<GID>212</GID>
<name>OUT_0</name></connection>
<intersection>-59.5 11</intersection>
<intersection>-50.5 12</intersection>
<intersection>-41.5 13</intersection>
<intersection>-32.5 14</intersection>
<intersection>-23.5 15</intersection>
<intersection>-14.5 4</intersection>
<intersection>-5.5 5</intersection>
<intersection>3.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15.5,3.5,41,3.5</points>
<connection>
<GID>192</GID>
<name>IN_0</name></connection>
<intersection>15.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>15.5,-14.5,41,-14.5</points>
<connection>
<GID>196</GID>
<name>IN_0</name></connection>
<intersection>15.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>15.5,-5.5,41,-5.5</points>
<connection>
<GID>194</GID>
<name>IN_0</name></connection>
<intersection>15.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>15.5,-59.5,41,-59.5</points>
<connection>
<GID>206</GID>
<name>IN_0</name></connection>
<intersection>15.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>15.5,-50.5,41,-50.5</points>
<connection>
<GID>204</GID>
<name>IN_0</name></connection>
<intersection>15.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>15.5,-41.5,41,-41.5</points>
<connection>
<GID>202</GID>
<name>IN_0</name></connection>
<intersection>15.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>15.5,-32.5,41,-32.5</points>
<connection>
<GID>200</GID>
<name>IN_0</name></connection>
<intersection>15.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>15.5,-23.5,41,-23.5</points>
<connection>
<GID>198</GID>
<name>IN_0</name></connection>
<intersection>15.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-10.5,-65.5,-10.5,5.5</points>
<connection>
<GID>214</GID>
<name>OUT_0</name></connection>
<intersection>-65.5 3</intersection>
<intersection>-47.5 8</intersection>
<intersection>-29.5 6</intersection>
<intersection>-11.5 4</intersection>
<intersection>5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-10.5,5,-9,5</points>
<connection>
<GID>216</GID>
<name>IN_0</name></connection>
<intersection>-10.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-10.5,-65.5,41,-65.5</points>
<connection>
<GID>206</GID>
<name>IN_3</name></connection>
<intersection>-10.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-10.5,-11.5,41,-11.5</points>
<connection>
<GID>194</GID>
<name>IN_3</name></connection>
<intersection>-10.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-10.5,-29.5,41,-29.5</points>
<connection>
<GID>198</GID>
<name>IN_3</name></connection>
<intersection>-10.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-10.5,-47.5,41,-47.5</points>
<connection>
<GID>202</GID>
<name>IN_3</name></connection>
<intersection>-10.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2,-63.5,-2,5.5</points>
<connection>
<GID>208</GID>
<name>OUT_0</name></connection>
<intersection>-63.5 9</intersection>
<intersection>-56.5 3</intersection>
<intersection>-27.5 7</intersection>
<intersection>-18.5 5</intersection>
<intersection>5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2,5,0,5</points>
<connection>
<GID>218</GID>
<name>IN_0</name></connection>
<intersection>-2 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-2,-56.5,41,-56.5</points>
<connection>
<GID>204</GID>
<name>IN_3</name></connection>
<intersection>-2 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-2,-18.5,41,-18.5</points>
<connection>
<GID>196</GID>
<name>IN_2</name></connection>
<intersection>-2 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-2,-27.5,41,-27.5</points>
<connection>
<GID>198</GID>
<name>IN_2</name></connection>
<intersection>-2 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-2,-63.5,41,-63.5</points>
<connection>
<GID>206</GID>
<name>IN_2</name></connection>
<intersection>-2 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6.5,-61.5,6.5,5.5</points>
<connection>
<GID>210</GID>
<name>OUT_0</name></connection>
<intersection>-61.5 9</intersection>
<intersection>-54.5 7</intersection>
<intersection>-43.5 5</intersection>
<intersection>-34.5 3</intersection>
<intersection>5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6.5,5,9,5</points>
<connection>
<GID>220</GID>
<name>IN_0</name></connection>
<intersection>6.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>6.5,-34.5,41,-34.5</points>
<connection>
<GID>200</GID>
<name>IN_1</name></connection>
<intersection>6.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>6.5,-43.5,41,-43.5</points>
<connection>
<GID>202</GID>
<name>IN_1</name></connection>
<intersection>6.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>6.5,-54.5,41,-54.5</points>
<connection>
<GID>204</GID>
<name>IN_2</name></connection>
<intersection>6.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>6.5,-61.5,41,-61.5</points>
<connection>
<GID>206</GID>
<name>IN_1</name></connection>
<intersection>6.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5,-52.5,-5,5</points>
<connection>
<GID>216</GID>
<name>OUT_0</name></connection>
<intersection>-52.5 7</intersection>
<intersection>-38.5 5</intersection>
<intersection>-20.5 3</intersection>
<intersection>-2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-5,-2.5,41,-2.5</points>
<connection>
<GID>192</GID>
<name>IN_3</name></connection>
<intersection>-5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-5,-20.5,41,-20.5</points>
<connection>
<GID>196</GID>
<name>IN_3</name></connection>
<intersection>-5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-5,-38.5,41,-38.5</points>
<connection>
<GID>200</GID>
<name>IN_3</name></connection>
<intersection>-5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-5,-52.5,41,-52.5</points>
<connection>
<GID>204</GID>
<name>IN_1</name></connection>
<intersection>-5 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4,-45.5,4,5</points>
<connection>
<GID>218</GID>
<name>OUT_0</name></connection>
<intersection>-45.5 5</intersection>
<intersection>-36.5 7</intersection>
<intersection>-9.5 3</intersection>
<intersection>-0.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>4,-0.5,41,-0.5</points>
<connection>
<GID>192</GID>
<name>IN_2</name></connection>
<intersection>4 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>4,-9.5,41,-9.5</points>
<connection>
<GID>194</GID>
<name>IN_2</name></connection>
<intersection>4 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>4,-45.5,41,-45.5</points>
<connection>
<GID>202</GID>
<name>IN_2</name></connection>
<intersection>4 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>4,-36.5,41,-36.5</points>
<connection>
<GID>200</GID>
<name>IN_2</name></connection>
<intersection>4 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-25.5,13,5</points>
<connection>
<GID>220</GID>
<name>OUT_0</name></connection>
<intersection>-25.5 5</intersection>
<intersection>-16.5 6</intersection>
<intersection>-7.5 7</intersection>
<intersection>1.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13,1.5,41,1.5</points>
<connection>
<GID>192</GID>
<name>IN_1</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>13,-25.5,41,-25.5</points>
<connection>
<GID>198</GID>
<name>IN_1</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>13,-16.5,41,-16.5</points>
<connection>
<GID>196</GID>
<name>IN_1</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>13,-7.5,41,-7.5</points>
<connection>
<GID>194</GID>
<name>IN_1</name></connection>
<intersection>13 0</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,0.5,47,0.5</points>
<connection>
<GID>224</GID>
<name>N_in0</name></connection>
<connection>
<GID>192</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-8.5,47,-8.5</points>
<connection>
<GID>226</GID>
<name>N_in0</name></connection>
<connection>
<GID>194</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-17.5,47,-17.5</points>
<connection>
<GID>228</GID>
<name>N_in0</name></connection>
<connection>
<GID>196</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-26.5,47,-26.5</points>
<connection>
<GID>230</GID>
<name>N_in0</name></connection>
<connection>
<GID>198</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-35.5,47,-35.5</points>
<connection>
<GID>232</GID>
<name>N_in0</name></connection>
<connection>
<GID>200</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-44.5,47,-44.5</points>
<connection>
<GID>234</GID>
<name>N_in0</name></connection>
<connection>
<GID>202</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-53.5,47,-53.5</points>
<connection>
<GID>236</GID>
<name>N_in0</name></connection>
<connection>
<GID>204</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-62.5,47,-62.5</points>
<connection>
<GID>238</GID>
<name>N_in0</name></connection>
<connection>
<GID>206</GID>
<name>OUT</name></connection></vsegment></shape></wire></page 3>
<page 4>
<PageViewport>-37.4,5.23333,125.8,-75.4333</PageViewport>
<gate>
<ID>386</ID>
<type>AA_TOGGLE</type>
<position>9,-155</position>
<output>
<ID>OUT_0</ID>129 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>388</ID>
<type>AA_TOGGLE</type>
<position>9,-160</position>
<output>
<ID>OUT_0</ID>130 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>390</ID>
<type>AA_TOGGLE</type>
<position>9,-164</position>
<output>
<ID>OUT_0</ID>131 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>392</ID>
<type>AA_TOGGLE</type>
<position>9,-170</position>
<output>
<ID>OUT_0</ID>132 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>394</ID>
<type>AA_LABEL</type>
<position>-0.5,-109.5</position>
<gparam>LABEL_TEXT 2*4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>396</ID>
<type>AA_LABEL</type>
<position>54.5,-107.5</position>
<gparam>LABEL_TEXT 3*8</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>398</ID>
<type>AA_LABEL</type>
<position>23,-137</position>
<gparam>LABEL_TEXT 4*16 DECODER </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>249</ID>
<type>AA_TOGGLE</type>
<position>22,-6</position>
<output>
<ID>OUT_0</ID>76 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>251</ID>
<type>AA_TOGGLE</type>
<position>30.5,-6</position>
<output>
<ID>OUT_0</ID>74 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>253</ID>
<type>AA_TOGGLE</type>
<position>39,-6</position>
<output>
<ID>OUT_0</ID>75 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>255</ID>
<type>AA_TOGGLE</type>
<position>46,-6</position>
<output>
<ID>OUT_0</ID>73 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>257</ID>
<type>AA_TOGGLE</type>
<position>53.5,-6</position>
<output>
<ID>OUT_0</ID>72 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>259</ID>
<type>AA_TOGGLE</type>
<position>61,-6</position>
<output>
<ID>OUT_0</ID>71 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>261</ID>
<type>AA_TOGGLE</type>
<position>68.5,-6</position>
<output>
<ID>OUT_0</ID>70 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>267</ID>
<type>AE_OR4</type>
<position>78.5,-17.5</position>
<input>
<ID>IN_0</ID>70 </input>
<input>
<ID>IN_1</ID>71 </input>
<input>
<ID>IN_2</ID>72 </input>
<input>
<ID>IN_3</ID>73 </input>
<output>
<ID>OUT</ID>77 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>269</ID>
<type>AE_OR4</type>
<position>78.5,-29.5</position>
<input>
<ID>IN_0</ID>74 </input>
<input>
<ID>IN_1</ID>75 </input>
<input>
<ID>IN_2</ID>71 </input>
<input>
<ID>IN_3</ID>70 </input>
<output>
<ID>OUT</ID>78 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>271</ID>
<type>AE_OR4</type>
<position>78.5,-41</position>
<input>
<ID>IN_0</ID>76 </input>
<input>
<ID>IN_1</ID>75 </input>
<input>
<ID>IN_2</ID>72 </input>
<input>
<ID>IN_3</ID>70 </input>
<output>
<ID>OUT</ID>79 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>273</ID>
<type>AA_TOGGLE</type>
<position>14.5,-6</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>275</ID>
<type>GA_LED</type>
<position>83.5,-17.5</position>
<input>
<ID>N_in0</ID>77 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>277</ID>
<type>GA_LED</type>
<position>83.5,-29.5</position>
<input>
<ID>N_in0</ID>78 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>279</ID>
<type>GA_LED</type>
<position>83.5,-41</position>
<input>
<ID>N_in0</ID>79 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>281</ID>
<type>AA_LABEL</type>
<position>14,-1.5</position>
<gparam>LABEL_TEXT OCTAL TO BINARY 8*3 DECODER </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>283</ID>
<type>AA_LABEL</type>
<position>14.5,-9.5</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>284</ID>
<type>AA_LABEL</type>
<position>23.5,-9</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>285</ID>
<type>AA_LABEL</type>
<position>32.5,-9</position>
<gparam>LABEL_TEXT D2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>286</ID>
<type>AA_LABEL</type>
<position>41,-9</position>
<gparam>LABEL_TEXT D3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>287</ID>
<type>AA_LABEL</type>
<position>47.5,-9.5</position>
<gparam>LABEL_TEXT D4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>288</ID>
<type>AA_LABEL</type>
<position>55.5,-9.5</position>
<gparam>LABEL_TEXT D5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>289</ID>
<type>AA_LABEL</type>
<position>62.5,-9.5</position>
<gparam>LABEL_TEXT D6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>290</ID>
<type>AA_LABEL</type>
<position>70.5,-9.5</position>
<gparam>LABEL_TEXT D7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>292</ID>
<type>AA_LABEL</type>
<position>90,-17</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>293</ID>
<type>AA_LABEL</type>
<position>89.5,-29</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>294</ID>
<type>AA_LABEL</type>
<position>89.5,-40.5</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>296</ID>
<type>AA_TOGGLE</type>
<position>25.5,-65</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>298</ID>
<type>AA_TOGGLE</type>
<position>39,-65</position>
<output>
<ID>OUT_0</ID>82 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>300</ID>
<type>AA_TOGGLE</type>
<position>50.5,-65</position>
<output>
<ID>OUT_0</ID>80 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>302</ID>
<type>AA_TOGGLE</type>
<position>64.5,-65</position>
<output>
<ID>OUT_0</ID>81 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>304</ID>
<type>AE_OR2</type>
<position>78.5,-75.5</position>
<input>
<ID>IN_0</ID>80 </input>
<input>
<ID>IN_1</ID>81 </input>
<output>
<ID>OUT</ID>83 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>308</ID>
<type>AE_OR2</type>
<position>79,-90.5</position>
<input>
<ID>IN_0</ID>82 </input>
<input>
<ID>IN_1</ID>81 </input>
<output>
<ID>OUT</ID>84 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>310</ID>
<type>GA_LED</type>
<position>82.5,-75.5</position>
<input>
<ID>N_in0</ID>83 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>312</ID>
<type>GA_LED</type>
<position>83,-90.5</position>
<input>
<ID>N_in0</ID>84 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>313</ID>
<type>AA_LABEL</type>
<position>26,-62</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>314</ID>
<type>AA_LABEL</type>
<position>39,-61.5</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>315</ID>
<type>AA_LABEL</type>
<position>50.5,-61</position>
<gparam>LABEL_TEXT D2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>316</ID>
<type>AA_LABEL</type>
<position>64,-60.5</position>
<gparam>LABEL_TEXT D3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>317</ID>
<type>AA_LABEL</type>
<position>87.5,-75</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>318</ID>
<type>AA_LABEL</type>
<position>88.5,-89.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>320</ID>
<type>AA_LABEL</type>
<position>22.5,-56</position>
<gparam>LABEL_TEXT 4*2 DECODER</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>322</ID>
<type>BA_DECODER_2x4</type>
<position>9,-120.5</position>
<input>
<ID>ENABLE</ID>85 </input>
<input>
<ID>IN_0</ID>87 </input>
<input>
<ID>IN_1</ID>86 </input>
<output>
<ID>OUT_0</ID>99 </output>
<output>
<ID>OUT_1</ID>98 </output>
<output>
<ID>OUT_2</ID>97 </output>
<output>
<ID>OUT_3</ID>96 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>324</ID>
<type>BE_DECODER_3x8</type>
<position>60,-120.5</position>
<input>
<ID>ENABLE</ID>88 </input>
<input>
<ID>IN_0</ID>91 </input>
<input>
<ID>IN_1</ID>90 </input>
<input>
<ID>IN_2</ID>89 </input>
<output>
<ID>OUT_0</ID>106 </output>
<output>
<ID>OUT_1</ID>107 </output>
<output>
<ID>OUT_2</ID>108 </output>
<output>
<ID>OUT_3</ID>105 </output>
<output>
<ID>OUT_4</ID>104 </output>
<output>
<ID>OUT_5</ID>103 </output>
<output>
<ID>OUT_6</ID>102 </output>
<output>
<ID>OUT_7</ID>100 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>326</ID>
<type>AA_TOGGLE</type>
<position>-0.5,-117</position>
<output>
<ID>OUT_0</ID>85 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>328</ID>
<type>AA_TOGGLE</type>
<position>-1,-120.5</position>
<output>
<ID>OUT_0</ID>86 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>330</ID>
<type>AA_TOGGLE</type>
<position>-1,-125</position>
<output>
<ID>OUT_0</ID>87 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>332</ID>
<type>AA_TOGGLE</type>
<position>53,-115</position>
<output>
<ID>OUT_0</ID>88 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>334</ID>
<type>AA_TOGGLE</type>
<position>53,-119</position>
<output>
<ID>OUT_0</ID>89 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>336</ID>
<type>AA_TOGGLE</type>
<position>52,-122.5</position>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>338</ID>
<type>AA_TOGGLE</type>
<position>52.5,-126</position>
<output>
<ID>OUT_0</ID>91 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>340</ID>
<type>GA_LED</type>
<position>19,-117</position>
<input>
<ID>N_in0</ID>96 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>344</ID>
<type>BI_DECODER_4x16</type>
<position>23.5,-155.5</position>
<input>
<ID>ENABLE</ID>128 </input>
<input>
<ID>IN_0</ID>132 </input>
<input>
<ID>IN_1</ID>131 </input>
<input>
<ID>IN_2</ID>130 </input>
<input>
<ID>IN_3</ID>129 </input>
<output>
<ID>OUT_0</ID>127 </output>
<output>
<ID>OUT_1</ID>112 </output>
<output>
<ID>OUT_10</ID>117 </output>
<output>
<ID>OUT_11</ID>116 </output>
<output>
<ID>OUT_12</ID>115 </output>
<output>
<ID>OUT_13</ID>109 </output>
<output>
<ID>OUT_14</ID>114 </output>
<output>
<ID>OUT_15</ID>113 </output>
<output>
<ID>OUT_2</ID>126 </output>
<output>
<ID>OUT_3</ID>125 </output>
<output>
<ID>OUT_4</ID>124 </output>
<output>
<ID>OUT_5</ID>111 </output>
<output>
<ID>OUT_6</ID>123 </output>
<output>
<ID>OUT_7</ID>122 </output>
<output>
<ID>OUT_8</ID>118 </output>
<output>
<ID>OUT_9</ID>110 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>346</ID>
<type>GA_LED</type>
<position>18,-120.5</position>
<input>
<ID>N_in0</ID>97 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>348</ID>
<type>GA_LED</type>
<position>18.5,-124</position>
<input>
<ID>N_in0</ID>98 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>350</ID>
<type>GA_LED</type>
<position>17.5,-128</position>
<input>
<ID>N_in0</ID>99 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>352</ID>
<type>GA_LED</type>
<position>72.5,-118.5</position>
<input>
<ID>N_in0</ID>103 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>354</ID>
<type>GA_LED</type>
<position>72.5,-121</position>
<input>
<ID>N_in0</ID>104 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>356</ID>
<type>GA_LED</type>
<position>69,-116</position>
<input>
<ID>N_in2</ID>102 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>358</ID>
<type>GA_LED</type>
<position>72.5,-124.5</position>
<input>
<ID>N_in0</ID>105 </input>
<input>
<ID>N_in3</ID>105 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>360</ID>
<type>GA_LED</type>
<position>65.5,-114.5</position>
<input>
<ID>N_in2</ID>100 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>362</ID>
<type>GA_LED</type>
<position>72.5,-127</position>
<input>
<ID>N_in0</ID>108 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>364</ID>
<type>GA_LED</type>
<position>68.5,-129.5</position>
<input>
<ID>N_in3</ID>107 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>366</ID>
<type>GA_LED</type>
<position>63,-130.5</position>
<input>
<ID>N_in3</ID>106 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>367</ID>
<type>GA_LED</type>
<position>44,-137.5</position>
<input>
<ID>N_in0</ID>113 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>368</ID>
<type>GA_LED</type>
<position>44,-140</position>
<input>
<ID>N_in0</ID>114 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>369</ID>
<type>GA_LED</type>
<position>44,-143.5</position>
<input>
<ID>N_in0</ID>109 </input>
<input>
<ID>N_in3</ID>109 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>370</ID>
<type>GA_LED</type>
<position>44,-146</position>
<input>
<ID>N_in0</ID>115 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>371</ID>
<type>GA_LED</type>
<position>44,-148.5</position>
<input>
<ID>N_in0</ID>116 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>372</ID>
<type>GA_LED</type>
<position>44,-151</position>
<input>
<ID>N_in0</ID>117 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>373</ID>
<type>GA_LED</type>
<position>44,-154.5</position>
<input>
<ID>N_in0</ID>110 </input>
<input>
<ID>N_in3</ID>110 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>374</ID>
<type>GA_LED</type>
<position>44,-157</position>
<input>
<ID>N_in0</ID>118 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>375</ID>
<type>GA_LED</type>
<position>44,-159.5</position>
<input>
<ID>N_in0</ID>122 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>376</ID>
<type>GA_LED</type>
<position>44,-162</position>
<input>
<ID>N_in0</ID>123 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>377</ID>
<type>GA_LED</type>
<position>44,-165.5</position>
<input>
<ID>N_in0</ID>111 </input>
<input>
<ID>N_in3</ID>111 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>378</ID>
<type>GA_LED</type>
<position>44,-168</position>
<input>
<ID>N_in0</ID>124 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>379</ID>
<type>GA_LED</type>
<position>44,-171.5</position>
<input>
<ID>N_in0</ID>125 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>380</ID>
<type>GA_LED</type>
<position>44,-174</position>
<input>
<ID>N_in0</ID>126 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>381</ID>
<type>GA_LED</type>
<position>44,-177.5</position>
<input>
<ID>N_in0</ID>112 </input>
<input>
<ID>N_in3</ID>112 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>382</ID>
<type>GA_LED</type>
<position>44,-180</position>
<input>
<ID>N_in0</ID>127 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>384</ID>
<type>AA_TOGGLE</type>
<position>18.5,-148</position>
<output>
<ID>OUT_0</ID>128 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-44,68.5,-8</points>
<connection>
<GID>261</GID>
<name>OUT_0</name></connection>
<intersection>-44 5</intersection>
<intersection>-32.5 3</intersection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68.5,-14.5,75.5,-14.5</points>
<connection>
<GID>267</GID>
<name>IN_0</name></connection>
<intersection>68.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>68.5,-32.5,75.5,-32.5</points>
<connection>
<GID>269</GID>
<name>IN_3</name></connection>
<intersection>68.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>68.5,-44,75.5,-44</points>
<connection>
<GID>271</GID>
<name>IN_3</name></connection>
<intersection>68.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,-30.5,61,-8</points>
<connection>
<GID>259</GID>
<name>OUT_0</name></connection>
<intersection>-30.5 3</intersection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61,-16.5,75.5,-16.5</points>
<connection>
<GID>267</GID>
<name>IN_1</name></connection>
<intersection>61 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>61,-30.5,75.5,-30.5</points>
<connection>
<GID>269</GID>
<name>IN_2</name></connection>
<intersection>61 0</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,-42,53.5,-8</points>
<connection>
<GID>257</GID>
<name>OUT_0</name></connection>
<intersection>-42 3</intersection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53.5,-18.5,75.5,-18.5</points>
<connection>
<GID>267</GID>
<name>IN_2</name></connection>
<intersection>53.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>53.5,-42,75.5,-42</points>
<connection>
<GID>271</GID>
<name>IN_2</name></connection>
<intersection>53.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-20.5,46,-8</points>
<connection>
<GID>255</GID>
<name>OUT_0</name></connection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-20.5,75.5,-20.5</points>
<connection>
<GID>267</GID>
<name>IN_3</name></connection>
<intersection>46 0</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-26.5,30.5,-8</points>
<connection>
<GID>251</GID>
<name>OUT_0</name></connection>
<intersection>-26.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-26.5,75.5,-26.5</points>
<connection>
<GID>269</GID>
<name>IN_0</name></connection>
<intersection>30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-40,39,-8</points>
<connection>
<GID>253</GID>
<name>OUT_0</name></connection>
<intersection>-40 3</intersection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-28.5,75.5,-28.5</points>
<connection>
<GID>269</GID>
<name>IN_1</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>39,-40,75.5,-40</points>
<connection>
<GID>271</GID>
<name>IN_1</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-38,22,-8</points>
<connection>
<GID>249</GID>
<name>OUT_0</name></connection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22,-38,75.5,-38</points>
<connection>
<GID>271</GID>
<name>IN_0</name></connection>
<intersection>22 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82.5,-17.5,82.5,-17.5</points>
<connection>
<GID>267</GID>
<name>OUT</name></connection>
<connection>
<GID>275</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82.5,-29.5,82.5,-29.5</points>
<connection>
<GID>269</GID>
<name>OUT</name></connection>
<connection>
<GID>277</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82.5,-41,82.5,-41</points>
<connection>
<GID>271</GID>
<name>OUT</name></connection>
<connection>
<GID>279</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-74.5,50.5,-67</points>
<connection>
<GID>300</GID>
<name>OUT_0</name></connection>
<intersection>-74.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-74.5,75.5,-74.5</points>
<connection>
<GID>304</GID>
<name>IN_0</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64.5,-91.5,64.5,-67</points>
<connection>
<GID>302</GID>
<name>OUT_0</name></connection>
<intersection>-91.5 3</intersection>
<intersection>-76.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64.5,-76.5,75.5,-76.5</points>
<connection>
<GID>304</GID>
<name>IN_1</name></connection>
<intersection>64.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>64.5,-91.5,76,-91.5</points>
<connection>
<GID>308</GID>
<name>IN_1</name></connection>
<intersection>64.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-89.5,39,-67</points>
<connection>
<GID>298</GID>
<name>OUT_0</name></connection>
<intersection>-89.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-89.5,76,-89.5</points>
<connection>
<GID>308</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81.5,-75.5,81.5,-75.5</points>
<connection>
<GID>304</GID>
<name>OUT</name></connection>
<connection>
<GID>310</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82,-90.5,82,-90.5</points>
<connection>
<GID>308</GID>
<name>OUT</name></connection>
<connection>
<GID>312</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3.5,-119,3.5,-117</points>
<intersection>-119 2</intersection>
<intersection>-117 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1.5,-117,3.5,-117</points>
<connection>
<GID>326</GID>
<name>OUT_0</name></connection>
<intersection>3.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>3.5,-119,6,-119</points>
<connection>
<GID>322</GID>
<name>ENABLE</name></connection>
<intersection>3.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3.5,-121,3.5,-120.5</points>
<intersection>-121 2</intersection>
<intersection>-120.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1,-120.5,3.5,-120.5</points>
<connection>
<GID>328</GID>
<name>OUT_0</name></connection>
<intersection>3.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>3.5,-121,6,-121</points>
<connection>
<GID>322</GID>
<name>IN_1</name></connection>
<intersection>3.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3.5,-125,3.5,-122</points>
<intersection>-125 1</intersection>
<intersection>-122 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1,-125,3.5,-125</points>
<connection>
<GID>330</GID>
<name>OUT_0</name></connection>
<intersection>3.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>3.5,-122,6,-122</points>
<connection>
<GID>322</GID>
<name>IN_0</name></connection>
<intersection>3.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-117,56,-115</points>
<intersection>-117 2</intersection>
<intersection>-115 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55,-115,56,-115</points>
<connection>
<GID>332</GID>
<name>OUT_0</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56,-117,57,-117</points>
<connection>
<GID>324</GID>
<name>ENABLE</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-122,56,-119</points>
<intersection>-122 2</intersection>
<intersection>-119 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55,-119,56,-119</points>
<connection>
<GID>334</GID>
<name>OUT_0</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56,-122,57,-122</points>
<connection>
<GID>324</GID>
<name>IN_2</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54,-123,57,-123</points>
<connection>
<GID>324</GID>
<name>IN_1</name></connection>
<intersection>54 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>54,-123,54,-122.5</points>
<connection>
<GID>336</GID>
<name>OUT_0</name></connection>
<intersection>-123 1</intersection></vsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-126,56,-124</points>
<intersection>-126 1</intersection>
<intersection>-124 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,-126,56,-126</points>
<connection>
<GID>338</GID>
<name>OUT_0</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56,-124,57,-124</points>
<connection>
<GID>324</GID>
<name>IN_0</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15,-119,15,-117</points>
<intersection>-119 2</intersection>
<intersection>-117 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,-117,18,-117</points>
<connection>
<GID>340</GID>
<name>N_in0</name></connection>
<intersection>15 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>12,-119,15,-119</points>
<connection>
<GID>322</GID>
<name>OUT_3</name></connection>
<intersection>15 0</intersection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-120.5,14.5,-120</points>
<intersection>-120.5 1</intersection>
<intersection>-120 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14.5,-120.5,17,-120.5</points>
<connection>
<GID>346</GID>
<name>N_in0</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>12,-120,14.5,-120</points>
<connection>
<GID>322</GID>
<name>OUT_2</name></connection>
<intersection>14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-124,14.5,-121</points>
<intersection>-124 1</intersection>
<intersection>-121 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14.5,-124,17.5,-124</points>
<connection>
<GID>348</GID>
<name>N_in0</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>12,-121,14.5,-121</points>
<connection>
<GID>322</GID>
<name>OUT_1</name></connection>
<intersection>14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14,-128,14,-122</points>
<intersection>-128 1</intersection>
<intersection>-122 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14,-128,16.5,-128</points>
<connection>
<GID>350</GID>
<name>N_in0</name></connection>
<intersection>14 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>12,-122,14,-122</points>
<connection>
<GID>322</GID>
<name>OUT_0</name></connection>
<intersection>14 0</intersection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,-117,65.5,-115.5</points>
<connection>
<GID>360</GID>
<name>N_in2</name></connection>
<intersection>-117 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63,-117,65.5,-117</points>
<connection>
<GID>324</GID>
<name>OUT_7</name></connection>
<intersection>65.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,-118,69,-117</points>
<connection>
<GID>356</GID>
<name>N_in2</name></connection>
<intersection>-118 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63,-118,69,-118</points>
<connection>
<GID>324</GID>
<name>OUT_6</name></connection>
<intersection>69 0</intersection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67,-119,67,-118.5</points>
<intersection>-119 2</intersection>
<intersection>-118.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>67,-118.5,71.5,-118.5</points>
<connection>
<GID>352</GID>
<name>N_in0</name></connection>
<intersection>67 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63,-119,67,-119</points>
<connection>
<GID>324</GID>
<name>OUT_5</name></connection>
<intersection>67 0</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>63,-120.5,71.5,-120.5</points>
<intersection>63 3</intersection>
<intersection>71.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>63,-120.5,63,-120</points>
<connection>
<GID>324</GID>
<name>OUT_4</name></connection>
<intersection>-120.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>71.5,-121,71.5,-120.5</points>
<connection>
<GID>354</GID>
<name>N_in0</name></connection>
<intersection>-120.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67,-124.5,67,-121</points>
<intersection>-124.5 1</intersection>
<intersection>-121 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>67,-124.5,72.5,-124.5</points>
<connection>
<GID>358</GID>
<name>N_in0</name></connection>
<intersection>67 0</intersection>
<intersection>72.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63,-121,67,-121</points>
<connection>
<GID>324</GID>
<name>OUT_3</name></connection>
<intersection>67 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>72.5,-124.5,72.5,-123.5</points>
<connection>
<GID>358</GID>
<name>N_in3</name></connection>
<intersection>-124.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-129.5,63,-124</points>
<connection>
<GID>324</GID>
<name>OUT_0</name></connection>
<connection>
<GID>366</GID>
<name>N_in3</name></connection></vsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-128.5,68.5,-123</points>
<connection>
<GID>364</GID>
<name>N_in3</name></connection>
<intersection>-123 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63,-123,68.5,-123</points>
<connection>
<GID>324</GID>
<name>OUT_1</name></connection>
<intersection>68.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67,-127,67,-122</points>
<intersection>-127 1</intersection>
<intersection>-122 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>67,-127,71.5,-127</points>
<connection>
<GID>362</GID>
<name>N_in0</name></connection>
<intersection>67 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63,-122,67,-122</points>
<connection>
<GID>324</GID>
<name>OUT_2</name></connection>
<intersection>67 0</intersection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-143.5,44,-143.5</points>
<connection>
<GID>369</GID>
<name>N_in0</name></connection>
<intersection>34 4</intersection>
<intersection>44 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>44,-143.5,44,-142.5</points>
<connection>
<GID>369</GID>
<name>N_in3</name></connection>
<intersection>-143.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>34,-150,34,-143.5</points>
<intersection>-150 5</intersection>
<intersection>-143.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>26.5,-150,34,-150</points>
<connection>
<GID>344</GID>
<name>OUT_13</name></connection>
<intersection>34 4</intersection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-154,44,-154</points>
<connection>
<GID>344</GID>
<name>OUT_9</name></connection>
<intersection>43 4</intersection>
<intersection>44 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>44,-154,44,-153.5</points>
<connection>
<GID>373</GID>
<name>N_in3</name></connection>
<intersection>-154 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>43,-154.5,43,-154</points>
<connection>
<GID>373</GID>
<name>N_in0</name></connection>
<intersection>-154 1</intersection></vsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39.5,-160.5,44,-160.5</points>
<intersection>39.5 4</intersection>
<intersection>43 5</intersection>
<intersection>44 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>44,-164.5,44,-160.5</points>
<connection>
<GID>377</GID>
<name>N_in3</name></connection>
<intersection>-160.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>39.5,-160.5,39.5,-158</points>
<intersection>-160.5 1</intersection>
<intersection>-158 6</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>43,-165.5,43,-160.5</points>
<connection>
<GID>377</GID>
<name>N_in0</name></connection>
<intersection>-160.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>26.5,-158,39.5,-158</points>
<connection>
<GID>344</GID>
<name>OUT_5</name></connection>
<intersection>39.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-177.5,44,-177.5</points>
<connection>
<GID>381</GID>
<name>N_in0</name></connection>
<intersection>31.5 4</intersection>
<intersection>44 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>44,-177.5,44,-176.5</points>
<connection>
<GID>381</GID>
<name>N_in3</name></connection>
<intersection>-177.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>31.5,-177.5,31.5,-162</points>
<intersection>-177.5 1</intersection>
<intersection>-162 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>26.5,-162,31.5,-162</points>
<connection>
<GID>344</GID>
<name>OUT_1</name></connection>
<intersection>31.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-148,38.5,-137.5</points>
<intersection>-148 1</intersection>
<intersection>-137.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-148,38.5,-148</points>
<connection>
<GID>344</GID>
<name>OUT_15</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>38.5,-137.5,43,-137.5</points>
<connection>
<GID>367</GID>
<name>N_in0</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-149,38.5,-140</points>
<intersection>-149 1</intersection>
<intersection>-140 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-149,38.5,-149</points>
<connection>
<GID>344</GID>
<name>OUT_14</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>38.5,-140,43,-140</points>
<connection>
<GID>368</GID>
<name>N_in0</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-151,38.5,-146</points>
<intersection>-151 1</intersection>
<intersection>-146 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-151,38.5,-151</points>
<connection>
<GID>344</GID>
<name>OUT_12</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>38.5,-146,43,-146</points>
<connection>
<GID>370</GID>
<name>N_in0</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-152,38.5,-148.5</points>
<intersection>-152 1</intersection>
<intersection>-148.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-152,38.5,-152</points>
<connection>
<GID>344</GID>
<name>OUT_11</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>38.5,-148.5,43,-148.5</points>
<connection>
<GID>371</GID>
<name>N_in0</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-153,38.5,-151</points>
<intersection>-153 1</intersection>
<intersection>-151 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-153,38.5,-153</points>
<connection>
<GID>344</GID>
<name>OUT_10</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>38.5,-151,43,-151</points>
<connection>
<GID>372</GID>
<name>N_in0</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-157,38.5,-155</points>
<intersection>-157 2</intersection>
<intersection>-155 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-155,38.5,-155</points>
<connection>
<GID>344</GID>
<name>OUT_8</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>38.5,-157,43,-157</points>
<connection>
<GID>374</GID>
<name>N_in0</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-159.5,38.5,-156</points>
<intersection>-159.5 2</intersection>
<intersection>-156 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-156,38.5,-156</points>
<connection>
<GID>344</GID>
<name>OUT_7</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>38.5,-159.5,43,-159.5</points>
<connection>
<GID>375</GID>
<name>N_in0</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-162,38.5,-157</points>
<intersection>-162 1</intersection>
<intersection>-157 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38.5,-162,43,-162</points>
<connection>
<GID>376</GID>
<name>N_in0</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26.5,-157,38.5,-157</points>
<connection>
<GID>344</GID>
<name>OUT_6</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-168,38.5,-159</points>
<intersection>-168 1</intersection>
<intersection>-159 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38.5,-168,43,-168</points>
<connection>
<GID>378</GID>
<name>N_in0</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26.5,-159,38.5,-159</points>
<connection>
<GID>344</GID>
<name>OUT_4</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-171.5,38.5,-160</points>
<intersection>-171.5 1</intersection>
<intersection>-160 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38.5,-171.5,43,-171.5</points>
<connection>
<GID>379</GID>
<name>N_in0</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26.5,-160,38.5,-160</points>
<connection>
<GID>344</GID>
<name>OUT_3</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-174,38.5,-161</points>
<intersection>-174 1</intersection>
<intersection>-161 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38.5,-174,43,-174</points>
<connection>
<GID>380</GID>
<name>N_in0</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26.5,-161,38.5,-161</points>
<connection>
<GID>344</GID>
<name>OUT_2</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-180,28.5,-163</points>
<intersection>-180 1</intersection>
<intersection>-163 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28.5,-180,43,-180</points>
<connection>
<GID>382</GID>
<name>N_in0</name></connection>
<intersection>28.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26.5,-163,28.5,-163</points>
<connection>
<GID>344</GID>
<name>OUT_0</name></connection>
<intersection>28.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,-148,20.5,-148</points>
<connection>
<GID>344</GID>
<name>ENABLE</name></connection>
<connection>
<GID>384</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18.5,-160,18.5,-155</points>
<intersection>-160 1</intersection>
<intersection>-155 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18.5,-160,20.5,-160</points>
<connection>
<GID>344</GID>
<name>IN_3</name></connection>
<intersection>18.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11,-155,18.5,-155</points>
<connection>
<GID>386</GID>
<name>OUT_0</name></connection>
<intersection>18.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>11,-160,20.5,-160</points>
<connection>
<GID>388</GID>
<name>OUT_0</name></connection>
<intersection>20.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>20.5,-161,20.5,-160</points>
<connection>
<GID>344</GID>
<name>IN_2</name></connection>
<intersection>-160 1</intersection></vsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-164,18,-162</points>
<intersection>-164 2</intersection>
<intersection>-162 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-162,20.5,-162</points>
<connection>
<GID>344</GID>
<name>IN_1</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11,-164,18,-164</points>
<connection>
<GID>390</GID>
<name>OUT_0</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-170,18,-163</points>
<intersection>-170 2</intersection>
<intersection>-163 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-163,20.5,-163</points>
<connection>
<GID>344</GID>
<name>IN_0</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11,-170,18,-170</points>
<connection>
<GID>392</GID>
<name>OUT_0</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire></page 4>
<page 5>
<PageViewport>-7.10543e-015,-18,122.4,-78.5</PageViewport>
<gate>
<ID>400</ID>
<type>AI_XOR2</type>
<position>43,-14.5</position>
<input>
<ID>IN_0</ID>133 </input>
<input>
<ID>IN_1</ID>134 </input>
<output>
<ID>OUT</ID>137 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>402</ID>
<type>AI_XOR2</type>
<position>43,-21</position>
<input>
<ID>IN_0</ID>134 </input>
<input>
<ID>IN_1</ID>135 </input>
<output>
<ID>OUT</ID>138 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>404</ID>
<type>AI_XOR2</type>
<position>42.5,-27.5</position>
<input>
<ID>IN_0</ID>135 </input>
<input>
<ID>IN_1</ID>136 </input>
<output>
<ID>OUT</ID>139 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>406</ID>
<type>AA_TOGGLE</type>
<position>26,-7</position>
<output>
<ID>OUT_0</ID>133 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>408</ID>
<type>AA_TOGGLE</type>
<position>27,-14</position>
<output>
<ID>OUT_0</ID>134 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>410</ID>
<type>AA_TOGGLE</type>
<position>27.5,-21</position>
<output>
<ID>OUT_0</ID>135 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>412</ID>
<type>AA_TOGGLE</type>
<position>28,-28.5</position>
<output>
<ID>OUT_0</ID>136 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>414</ID>
<type>GA_LED</type>
<position>58,-7</position>
<input>
<ID>N_in0</ID>133 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>416</ID>
<type>GA_LED</type>
<position>58,-13</position>
<input>
<ID>N_in0</ID>137 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>418</ID>
<type>GA_LED</type>
<position>58,-20</position>
<input>
<ID>N_in0</ID>138 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>420</ID>
<type>GA_LED</type>
<position>58,-27</position>
<input>
<ID>N_in0</ID>139 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>422</ID>
<type>AA_LABEL</type>
<position>36.5,-2.5</position>
<gparam>LABEL_TEXT BINARY TO GRAY</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>424</ID>
<type>AA_LABEL</type>
<position>17,-6.5</position>
<gparam>LABEL_TEXT B4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>426</ID>
<type>AA_LABEL</type>
<position>65.5,-6.5</position>
<gparam>LABEL_TEXT G4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>427</ID>
<type>AA_LABEL</type>
<position>17.5,-14</position>
<gparam>LABEL_TEXT B3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>428</ID>
<type>AA_LABEL</type>
<position>20,-28.5</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>429</ID>
<type>AA_LABEL</type>
<position>18.5,-21</position>
<gparam>LABEL_TEXT B2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>430</ID>
<type>AA_LABEL</type>
<position>66,-13</position>
<gparam>LABEL_TEXT G3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>431</ID>
<type>AA_LABEL</type>
<position>65.5,-20</position>
<gparam>LABEL_TEXT G2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>432</ID>
<type>AA_LABEL</type>
<position>66,-26</position>
<gparam>LABEL_TEXT G1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>434</ID>
<type>AA_LABEL</type>
<position>35,-35.5</position>
<gparam>LABEL_TEXT GRAY  TO BINARY </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>436</ID>
<type>AA_TOGGLE</type>
<position>24.5,-44</position>
<output>
<ID>OUT_0</ID>149 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>438</ID>
<type>AA_TOGGLE</type>
<position>32,-44</position>
<output>
<ID>OUT_0</ID>145 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>440</ID>
<type>AA_TOGGLE</type>
<position>41,-44</position>
<output>
<ID>OUT_0</ID>144 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>442</ID>
<type>AA_TOGGLE</type>
<position>52.5,-44</position>
<output>
<ID>OUT_0</ID>143 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>444</ID>
<type>AI_XOR2</type>
<position>60.5,-52</position>
<input>
<ID>IN_0</ID>143 </input>
<input>
<ID>IN_1</ID>144 </input>
<output>
<ID>OUT</ID>140 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>448</ID>
<type>AI_XOR3</type>
<position>61,-60.5</position>
<input>
<ID>IN_0</ID>145 </input>
<input>
<ID>IN_1</ID>144 </input>
<input>
<ID>IN_2</ID>143 </input>
<output>
<ID>OUT</ID>141 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>452</ID>
<type>GA_LED</type>
<position>64.5,-52</position>
<input>
<ID>N_in0</ID>140 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>454</ID>
<type>GA_LED</type>
<position>65,-60.5</position>
<input>
<ID>N_in0</ID>141 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>456</ID>
<type>GA_LED</type>
<position>65,-70</position>
<input>
<ID>N_in0</ID>148 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>458</ID>
<type>GA_LED</type>
<position>64.5,-46.5</position>
<input>
<ID>N_in0</ID>143 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>462</ID>
<type>AI_XOR4</type>
<position>60,-70</position>
<input>
<ID>IN_0</ID>143 </input>
<input>
<ID>IN_1</ID>144 </input>
<input>
<ID>IN_2</ID>145 </input>
<input>
<ID>IN_3</ID>149 </input>
<output>
<ID>OUT</ID>148 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<wire>
<ID>133</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28,-7,57,-7</points>
<connection>
<GID>406</GID>
<name>OUT_0</name></connection>
<connection>
<GID>414</GID>
<name>N_in0</name></connection>
<intersection>36 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>36,-13.5,36,-7</points>
<intersection>-13.5 3</intersection>
<intersection>-7 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>36,-13.5,40,-13.5</points>
<connection>
<GID>400</GID>
<name>IN_0</name></connection>
<intersection>36 2</intersection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-20,34.5,-14</points>
<intersection>-20 4</intersection>
<intersection>-15.5 1</intersection>
<intersection>-14 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34.5,-15.5,40,-15.5</points>
<connection>
<GID>400</GID>
<name>IN_1</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-14,34.5,-14</points>
<connection>
<GID>408</GID>
<name>OUT_0</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>34.5,-20,40,-20</points>
<connection>
<GID>402</GID>
<name>IN_0</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-26.5,34.5,-21</points>
<intersection>-26.5 4</intersection>
<intersection>-22 2</intersection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29.5,-21,34.5,-21</points>
<connection>
<GID>410</GID>
<name>OUT_0</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34.5,-22,40,-22</points>
<connection>
<GID>402</GID>
<name>IN_1</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>34.5,-26.5,39.5,-26.5</points>
<connection>
<GID>404</GID>
<name>IN_0</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30,-28.5,39.5,-28.5</points>
<connection>
<GID>412</GID>
<name>OUT_0</name></connection>
<intersection>39.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>39.5,-28.5,39.5,-28.5</points>
<connection>
<GID>404</GID>
<name>IN_1</name></connection>
<intersection>-28.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,-14.5,51.5,-13</points>
<intersection>-14.5 2</intersection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51.5,-13,57,-13</points>
<connection>
<GID>416</GID>
<name>N_in0</name></connection>
<intersection>51.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>46,-14.5,51.5,-14.5</points>
<connection>
<GID>400</GID>
<name>OUT</name></connection>
<intersection>51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,-21,51.5,-20</points>
<intersection>-21 2</intersection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51.5,-20,57,-20</points>
<connection>
<GID>418</GID>
<name>N_in0</name></connection>
<intersection>51.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>46,-21,51.5,-21</points>
<connection>
<GID>402</GID>
<name>OUT</name></connection>
<intersection>51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-27.5,51,-27</points>
<intersection>-27.5 2</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51,-27,57,-27</points>
<connection>
<GID>420</GID>
<name>N_in0</name></connection>
<intersection>51 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45.5,-27.5,51,-27.5</points>
<connection>
<GID>404</GID>
<name>OUT</name></connection>
<intersection>51 0</intersection></hsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,-52,63.5,-52</points>
<connection>
<GID>452</GID>
<name>N_in0</name></connection>
<connection>
<GID>444</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,-60.5,64,-60.5</points>
<connection>
<GID>454</GID>
<name>N_in0</name></connection>
<connection>
<GID>448</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-67,52.5,-46</points>
<connection>
<GID>442</GID>
<name>OUT_0</name></connection>
<intersection>-67 8</intersection>
<intersection>-62.5 6</intersection>
<intersection>-51 4</intersection>
<intersection>-46.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52.5,-46.5,63.5,-46.5</points>
<connection>
<GID>458</GID>
<name>N_in0</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>52.5,-51,57.5,-51</points>
<connection>
<GID>444</GID>
<name>IN_0</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>52.5,-62.5,58,-62.5</points>
<connection>
<GID>448</GID>
<name>IN_2</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>52.5,-67,57,-67</points>
<connection>
<GID>462</GID>
<name>IN_0</name></connection>
<intersection>52.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41,-69,41,-46</points>
<connection>
<GID>440</GID>
<name>OUT_0</name></connection>
<intersection>-69 7</intersection>
<intersection>-60.5 3</intersection>
<intersection>-53 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41,-53,57.5,-53</points>
<connection>
<GID>444</GID>
<name>IN_1</name></connection>
<intersection>41 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>41,-60.5,58,-60.5</points>
<connection>
<GID>448</GID>
<name>IN_1</name></connection>
<intersection>41 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>41,-69,57,-69</points>
<connection>
<GID>462</GID>
<name>IN_1</name></connection>
<intersection>41 0</intersection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-71,32,-46</points>
<connection>
<GID>438</GID>
<name>OUT_0</name></connection>
<intersection>-71 5</intersection>
<intersection>-58.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,-58.5,58,-58.5</points>
<connection>
<GID>448</GID>
<name>IN_0</name></connection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>32,-71,57,-71</points>
<connection>
<GID>462</GID>
<name>IN_2</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,-70,64,-70</points>
<connection>
<GID>462</GID>
<name>OUT</name></connection>
<connection>
<GID>456</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-73,24.5,-46</points>
<connection>
<GID>436</GID>
<name>OUT_0</name></connection>
<intersection>-73 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-73,57,-73</points>
<connection>
<GID>462</GID>
<name>IN_3</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire></page 5>
<page 6>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 6>
<page 7>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 7>
<page 8>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 9></circuit>